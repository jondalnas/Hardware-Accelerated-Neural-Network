library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.types.all;
use IEEE.NUMERIC_STD.ALL;

entity nn is
    generic(
        num_in : positive;
        num_out : positive;
        num_feedback : positive;
        data_width : integer
    );
    Port (
        clk : in std_logic;
        rst : in std_logic;
        valid_in : in std_logic;
        valid_out : out std_logic;
        input : in array_type(num_in-1 downto 0);
        output : out array_type(num_out-1 downto 0)
     );
end nn;

architecture Behavioral of nn is
    signal feedback, next_feedback : array_type(num_feedback-1 downto 0)(data_width - 1 downto 0);
    signal was_valid, next_was_valid : std_logic;

    signal state, next_state : integer;

    signal Block386_o : array_type(783 downto 0)(data_width-1 downto 0);
    signal Block386_i_0 : array_type(783 downto 0)(data_width-1 downto 0);
    signal Block386_i_1 : array_type(0 downto 0)(data_width-1 downto 0);
    signal Block386_bc_i_1 : array_type(783 downto 0)(data_width-1 downto 0);
    signal Convolution28_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Convolution28_i_0 : array_type(783 downto 0)(data_width-1 downto 0);
    signal Convolution28_i_1 : array_type(199 downto 0)(data_width-1 downto 0);
    signal Plus30_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Plus30_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Plus30_i_1 : array_type(7 downto 0)(data_width-1 downto 0);
    signal Plus30_bc_i_1 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal ReLU32_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal ReLU32_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Pooling66_o : array_type(1567 downto 0)(data_width-1 downto 0);
    signal Pooling66_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Convolution110_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Convolution110_i_0 : array_type(1567 downto 0)(data_width-1 downto 0);
    signal Convolution110_i_1 : array_type(3199 downto 0)(data_width-1 downto 0);
    signal Plus112_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Plus112_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Plus112_i_1 : array_type(15 downto 0)(data_width-1 downto 0);
    signal Plus112_bc_i_1 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal ReLU114_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal ReLU114_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Pooling160_o : array_type(255 downto 0)(data_width-1 downto 0);
    signal Pooling160_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Times212_o : array_type(9 downto 0)(data_width-1 downto 0);
    signal Times212_i_0 : array_type(255 downto 0)(data_width-1 downto 0);
    signal Times212_i_1 : array_type(2559 downto 0)(data_width-1 downto 0);
    signal Plus214_o : array_type(9 downto 0)(data_width-1 downto 0);
    signal Plus214_i_0 : array_type(9 downto 0)(data_width-1 downto 0);
    signal Plus214_i_1 : array_type(9 downto 0)(data_width-1 downto 0);
    signal Block386_valid_in, Block386_valid_out, Convolution28_valid_in, Convolution28_valid_out, Plus30_valid_in, Plus30_valid_out, ReLU32_valid_in, ReLU32_valid_out, Pooling66_valid_in, Pooling66_valid_out, Convolution110_valid_in, Convolution110_valid_out, Plus112_valid_in, Plus112_valid_out, ReLU114_valid_in, ReLU114_valid_out, Pooling160_valid_in, Pooling160_valid_out, Times212_valid_in, Times212_valid_out, Plus214_valid_in, Plus214_valid_out : std_logic;
begin
    Block386 : entity work.div
        generic map (
            input_size => 784,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Block386_valid_in,
            valid_out => Block386_valid_out,
            a => Block386_i_0,
            b => Block386_bc_i_1,
            c => Block386_o
        );
    Block386_1_bc : entity work.broad
        generic map(
            input_size => 1,
            block_repeat => 1,
            element_repeat => 784,
            data_width => 16
        )
        port map(
            input => Block386_i_1,
            output => Block386_bc_i_1
        );
    Convolution28 : entity work.conv
        generic map (
            num_dimensions => 4,
            dimensions_x => (1, 1, 28, 28),
            x_size => 784,
            dimensions_w => (8, 1, 5, 5),
            w_size => 200,
            kernel_shape => (5, 5),
            kernel_size => 25,
            dilation => (1, 1),
            stride => (1, 1),
            data_width => 16,
            y_size => 6272
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Convolution28_valid_in,
            valid_out => Convolution28_valid_out,
            x => Convolution28_i_0,
            w => Convolution28_i_1,
            y => Convolution28_o
        );
    Plus30 : entity work.add
        generic map (
            input_size => 6272,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Plus30_valid_in,
            valid_out => Plus30_valid_out,
            a => Plus30_i_0,
            b => Plus30_bc_i_1,
            c => Plus30_o
        );
    Plus30_1_bc : entity work.broad
        generic map(
            input_size => 8,
            block_repeat => 1,
            element_repeat => 784,
            data_width => 16
        )
        port map(
            input => Plus30_i_1,
            output => Plus30_bc_i_1
        );
    ReLU32 : entity work.relu
        generic map (
            input_size => 6272,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => ReLU32_valid_in,
            valid_out => ReLU32_valid_out,
            x => ReLU32_i_0,
            y => ReLU32_o
        );
    Pooling66 : entity work.max_pool
        generic map (
            num_dimensions => 4,
            kernel_shape => (2, 2),
            pads => (0, 0, 0, 0),
            strides => (2, 2),
            in_dimensions => (1, 8, 28, 28),
            out_dimensions => (1, 8, 14, 14),
            input_size => 6272,
            output_size => 1568,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Pooling66_valid_in,
            valid_out => Pooling66_valid_out,
            x => Pooling66_i_0,
            y => Pooling66_o
        );
    Convolution110 : entity work.conv
        generic map (
            num_dimensions => 4,
            dimensions_x => (1, 8, 14, 14),
            x_size => 1568,
            dimensions_w => (16, 8, 5, 5),
            w_size => 3200,
            kernel_shape => (5, 5),
            kernel_size => 25,
            dilation => (1, 1),
            stride => (1, 1),
            data_width => 16,
            y_size => 3136
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Convolution110_valid_in,
            valid_out => Convolution110_valid_out,
            x => Convolution110_i_0,
            w => Convolution110_i_1,
            y => Convolution110_o
        );
    Plus112 : entity work.add
        generic map (
            input_size => 3136,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Plus112_valid_in,
            valid_out => Plus112_valid_out,
            a => Plus112_i_0,
            b => Plus112_bc_i_1,
            c => Plus112_o
        );
    Plus112_1_bc : entity work.broad
        generic map(
            input_size => 16,
            block_repeat => 1,
            element_repeat => 196,
            data_width => 16
        )
        port map(
            input => Plus112_i_1,
            output => Plus112_bc_i_1
        );
    ReLU114 : entity work.relu
        generic map (
            input_size => 3136,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => ReLU114_valid_in,
            valid_out => ReLU114_valid_out,
            x => ReLU114_i_0,
            y => ReLU114_o
        );
    Pooling160 : entity work.max_pool
        generic map (
            num_dimensions => 4,
            kernel_shape => (3, 3),
            pads => (0, 0, 0, 0),
            strides => (3, 3),
            in_dimensions => (1, 16, 14, 14),
            out_dimensions => (1, 16, 4, 4),
            input_size => 3136,
            output_size => 256,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Pooling160_valid_in,
            valid_out => Pooling160_valid_out,
            x => Pooling160_i_0,
            y => Pooling160_o
        );
    Times212 : entity work.mat_mul
        generic map (
            num_dimensions => 2,
            a_dim => (1, 256),
            b_dim => (256, 10),
            a_size => 256,
            b_size => 2560,
            y_size => 10,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Times212_valid_in,
            valid_out => Times212_valid_out,
            a => Times212_i_0,
            b => Times212_i_1,
            y => Times212_o
        );
    Plus214 : entity work.add
        generic map (
            input_size => 10,
            data_width => 16
        )
        port map (
            clk => clk,
            rst => rst,
            valid_in => Plus214_valid_in,
            valid_out => Plus214_valid_out,
            a => Plus214_i_0,
            b => Plus214_i_1,
            c => Plus214_o
        );

    Block386_i_1 <= (0 => "0111111111111111");
    Convolution28_i_1 <= ("1111111111010000", "1111111110111000", "1111111110010011", "1111111111010000", "1111111111110111", "1111111110000000", "1111111111001110", "1111111111100010", "1111111111011101", "0000000000000111", "0000000000100010", "0000000000001100", "0000000000100001", "0000000000110010", "1111111111100010", "0000000010010001", "0000000001010000", "0000000000110001", "0000000001100000", "0000000000101010", "0000000001010110", "0000000000111011", "0000000000010111", "1111111111011111", "1111111111111011", "1111111111110101", "0000000000100010", "0000000000010010", "0000000000101111", "0000000001011001", "1111111111011010", "1111111110100110", "1111111111010100", "0000000000011101", "0000000001000111", "1111111111101010", "1111111110110011", "1111111110001011", "0000000001001100", "0000000001101010", "1111111111000001", "1111111110010011", "1111111110011000", "0000000001111100", "0000000001011101", "1111111111001010", "1111111110001011", "1111111111001010", "0000000010001111", "0000000000011001", "0000000000111001", "0000000001111000", "0000000000111100", "0000000001001101", "0000000000001111", "1111111111100100", "0000000000100001", "0000000001011101", "0000000010101000", "0000000000111000", "1111111111001011", "1111111110101000", "1111111111000000", "0000000001011000", "0000000010001010", "1111111110011110", "1111111101101010", "1111111101000101", "1111111101110100", "0000000000101110", "0000000000100100", "0000000000001101", "1111111111010000", "1111111110101011", "1111111111010110", "0000000000111100", "0000000010101110", "0000000010100000", "0000000000111111", "0000000000000010", "1111111111111110", "0000000000001010", "0000000001000110", "0000000000100100", "1111111111100011", "1111111101110000", "1111111110000111", "1111111111111101", "0000000001101001", "1111111111110001", "1111111101110001", "1111111111000111", "1111111111011000", "0000000000110100", "0000000000010110", "1111111111010111", "1111111111000111", "0000000000000000", "1111111111100001", "1111111111001010", "0000000001010111", "0000000000110101", "0000000000000111", "0000000001011001", "0000000001010011", "0000000000101110", "1111111111111110", "0000000000111000", "0000000001011111", "0000000000011000", "0000000000111010", "0000000000001010", "0000000000011111", "1111111111111010", "1111111110011100", "0000000000101001", "0000000000101001", "1111111111110010", "1111111111001011", "1111111110000110", "1111111111001000", "1111111111101100", "1111111110101101", "1111111110101011", "1111111110110101", "1111111111110000", "1111111111011011", "1111111110100111", "1111111110101011", "1111111111001110", "1111111110001110", "1111111101100011", "1111111101110111", "1111111101001001", "1111111100000111", "1111111111000001", "1111111111010100", "1111111111011100", "1111111111101101", "1111111110001000", "0000000000111110", "0000000001010100", "0000000001100010", "0000000001101010", "0000000001010101", "0000000010110000", "0000000001011100", "0000000001000000", "0000000000011010", "1111111111111010", "0000000001001000", "1111111111111101", "1111111111110000", "1111111111000110", "1111111110011111", "0000000001010101", "0000000000111010", "1111111111010100", "1111111110011110", "1111111101101111", "0000000001011111", "0000000001011011", "1111111111011000", "1111111110101101", "1111111111011010", "0000000001100111", "0000000010000110", "1111111111111111", "1111111110111010", "1111111111100111", "0000000000001100", "0000000001101100", "0000000001111111", "0000000000110111", "1111111111110110", "1111111110110110", "1111111110000110", "1111111111001001", "0000000000111001", "0000000000001001", "1111111101100100", "1111111110110101", "0000000010010111", "0000000010001110", "1111111111011000", "1111111110001111", "0000000010001110", "0000000100000100", "0000000000001110", "1111111110000011", "0000000001000011", "0000000011000100", "1111111111110100", "1111111110000111", "1111111101101001", "0000000000100100", "1111111111110000", "1111111101111110", "1111111111000100", "1111111111111110");
    Plus30_i_1 <= ("1111111111100001", "0000000000000101", "1111111111011111", "1111111111110000", "1111111111111100", "0000000000010111", "1111111110010001", "1111111111010111");
    Convolution110_i_1 <= ("1111111111100011", "0000000000000011", "1111111111011100", "0000000000001101", "1111111111001011", "1111111111101000", "1111111111001011", "0000000000000000", "1111111111111111", "1111111111100110", "1111111111101000", "1111111111011100", "1111111111110000", "0000000000010001", "1111111110010010", "0000000000110010", "0000000000100001", "0000000000000011", "1111111111000001", "1111111110110010", "0000000000010001", "0000000000001111", "0000000000010000", "0000000000000001", "1111111111011011", "0000000000000000", "0000000000011000", "0000000000110100", "0000000001011101", "1111111111010111", "0000000000000010", "0000000000100001", "0000000000101010", "0000000000100101", "1111111111010001", "0000000000010111", "0000000000100100", "0000000000001010", "1111111111001100", "0000000000011000", "1111111111111010", "0000000000001000", "1111111111111101", "1111111110110010", "0000000000000001", "1111111111011110", "1111111111101010", "1111111111000011", "1111111111000110", "1111111111100010", "1111111111011100", "1111111111100111", "1111111111100100", "1111111111110000", "1111111111000000", "1111111111101111", "0000000000011101", "1111111111100100", "1111111111111110", "1111111111010100", "0000000000100011", "0000000000000110", "1111111111111101", "0000000000001011", "0000000000000100", "0000000000000010", "1111111111011000", "1111111111111010", "1111111111000001", "1111111111101010", "0000000000000011", "1111111111100111", "1111111110101111", "1111111110110000", "1111111111000110", "1111111111010001", "0000000000000011", "1111111111100100", "0000000000001000", "1111111111101010", "1111111111111100", "1111111111100000", "0000000000001010", "0000000000001011", "1111111111011100", "1111111111101101", "1111111111101010", "0000000000001101", "0000000000001000", "1111111111110011", "1111111111001010", "0000000000000001", "0000000000001111", "1111111111011011", "1111111110111000", "1111111111010111", "1111111111111001", "1111111111111000", "1111111110010110", "1111111110100111", "1111111111111100", "1111111111000100", "1111111111100101", "0000000000000011", "0000000001001011", "1111111111101011", "1111111110111001", "0000000000000000", "0000000001000000", "1111111111111100", "1111111111010011", "1111111111000011", "0000000000010100", "0000000001001101", "1111111111111000", "1111111111100111", "1111111111000011", "0000000000011010", "0000000000011110", "1111111111101011", "1111111111011110", "0000000000001101", "0000000000010000", "0000000000001100", "1111111110101100", "1111111111100010", "0000000000000010", "1111111111110010", "1111111111101001", "1111111110110010", "1111111111010000", "1111111111100001", "1111111111100001", "1111111111010010", "1111111111001110", "0000000000011100", "1111111111100000", "1111111110111111", "1111111111010011", "1111111111000010", "0000000000011110", "1111111111110100", "1111111111010010", "1111111111100101", "0000000000001100", "0000000000000011", "1111111111010010", "0000000000000111", "0000000000000011", "1111111111101011", "1111111111110000", "1111111111010110", "1111111111000101", "1111111111110000", "0000000000100011", "1111111111110110", "1111111110111110", "1111111111111100", "0000000000101101", "0000000000010101", "1111111111101010", "1111111111010100", "1111111111110110", "0000000001001111", "0000000000011100", "1111111111101010", "1111111111101001", "0000000000010010", "0000000001100000", "1111111111101111", "1111111111001100", "1111111111110011", "0000000000011000", "0000000001001100", "1111111111010111", "1111111111101111", "1111111111110100", "0000000000000101", "0000000000010000", "0000000000011010", "1111111111100100", "1111111111001111", "1111111111110010", "0000000000101101", "0000000000100110", "1111111111110001", "1111111111111010", "0000000000101100", "0000000000101100", "1111111111011111", "1111111111001110", "1111111111111011", "0000000000110111", "0000000000100100", "1111111110101111", "0000000000001001", "1111111111011011", "0000000000001000", "1111111111111010", "1111111110111101", "1111111111110111", "1111111111011001", "1111111111000010", "0000000000001001", "0000000000010100", "1111111111100011", "1111111111110000", "1111111111001110", "1111111111101001", "1111111111100111", "1111111111111001", "1111111111110011", "1111111111110110", "1111111111100111", "1111111111010000", "1111111111000110", "1111111111010111", "1111111111001001", "1111111111100000", "1111111111100011", "0000000000100011", "0000000000101111", "0000000000111100", "0000000000100111", "0000000000011101", "0000000000010100", "1111111111010101", "0000000000001101", "0000000001011111", "0000000000010100", "0000000000000101", "1111111111110101", "0000000000010111", "0000000001001010", "0000000000000000", "1111111111100110", "1111111111110000", "0000000000010101", "0000000000011001", "0000000000110110", "1111111111110110", "1111111111100001", "0000000000000010", "1111111111110011", "0000000000000101", "1111111111110011", "1111111111011101", "0000000000000001", "1111111111010100", "1111111111010001", "0000000000100101", "1111111111010001", "1111111111011010", "1111111111011100", "1111111111100001", "0000000000001111", "0000000000000000", "0000000000010001", "0000000000110010", "1111111111010100", "0000000000000001", "1111111111000101", "0000000000001110", "0000000001000010", "0000000000000000", "0000000000000111", "0000000000011001", "1111111111110000", "1111111111011000", "0000000000001101", "1111111111100111", "1111111111100101", "1111111111111010", "1111111111101011", "1111111111010001", "0000000000101111", "1111111111100111", "1111111111001010", "0000000000001100", "1111111111101101", "0000000000101101", "1111111111100100", "0000000000001101", "0000000000010110", "1111111111001011", "1111111111111010", "1111111111011010", "1111111111001101", "0000000000110000", "0000000000001010", "0000000000010101", "0000000000000001", "1111111111100101", "1111111111110101", "0000000000010010", "1111111111101111", "1111111111010110", "1111111111110100", "1111111111111100", "1111111110110101", "0000000000011110", "1111111111111101", "1111111111000000", "1111111111111100", "0000000000101110", "0000000000111110", "1111111111101000", "1111111110111001", "1111111111101101", "0000000000000101", "0000000000011111", "1111111111101100", "1111111111010000", "1111111111010011", "1111111111011100", "0000000000001010", "0000000000000001", "1111111111101000", "1111111111111011", "0000000000010101", "1111111111101010", "1111111111101001", "0000000000000000", "0000000000001010", "1111111111101000", "1111111111010010", "1111111110111011", "1111111111001011", "1111111111011101", "1111111111111000", "0000000000000001", "1111111111110101", "1111111111110001", "1111111111100110", "1111111111110111", "0000000000101010", "0000000000100100", "0000000000000100", "1111111111100100", "1111111111010001", "1111111111001110", "1111111111010010", "1111111111111110", "1111111111110000", "1111111111100111", "0000000000111000", "0000000000110101", "0000000000010100", "0000000000100010", "1111111111101101", "0000000000110111", "0000000001000111", "0000000000000010", "0000000000001000", "0000000001000011", "0000000000011001", "0000000000100100", "0000000000000111", "0000000000001101", "0000000000101101", "0000000000010101", "0000000000101011", "1111111111111010", "1111111111101101", "0000000000001110", "1111111111111111", "1111111111101101", "1111111111011001", "1111111111000101", "1111111111010111", "0000000000111011", "0000000000011011", "0000000000010110", "0000000000001100", "1111111111110001", "1111111111011111", "1111111111110110", "1111111111001010", "1111111111110110", "0000000001010000", "1111111110111010", "1111111111011100", "1111111111011101", "1111111111100110", "0000000000011001", "1111111111111100", "0000000000010001", "1111111111101000", "1111111111111000", "1111111111000100", "1111111111111000", "0000000000001010", "1111111111100011", "1111111111111010", "1111111111110111", "1111111111111001", "1111111111110100", "0000000000010100", "0000000000001111", "0000000000110110", "1111111111101010", "1111111111111001", "1111111111101001", "1111111111101100", "0000000000100101", "1111111111011100", "0000000000011010", "1111111111110100", "1111111111001011", "1111111111100000", "0000000000101000", "0000000000101011", "1111111111101010", "0000000000000111", "0000000000101000", "0000000000011110", "0000000000011111", "0000000000010010", "0000000000111011", "0000000000011000", "1111111110111111", "1111111111001101", "1111111111001110", "1111111111111001", "0000000000011011", "1111111111000000", "0000000001011100", "0000000001010011", "0000000000001011", "1111111111100001", "0000000001100110", "0000000001001010", "1111111111001001", "1111111111000001", "1111111111010101", "0000000000110100", "0000000000010010", "1111111110100101", "1111111110101011", "1111111110110001", "0000000000000111", "1111111111000100", "1111111110101110", "1111111111001110", "1111111111011000", "1111111111110111", "1111111111001111", "1111111111001011", "0000000000000111", "0000000000000001", "0000000000010101", "1111111111011100", "1111111111000100", "1111111111011000", "1111111111100011", "0000000000100101", "1111111111001110", "1111111110111000", "1111111111100110", "0000000000100111", "1111111111100000", "0000000000101010", "1111111111101010", "1111111111100001", "1111111111111101", "1111111111100011", "1111111111101011", "0000000000001100", "0000000000010010", "0000000000011101", "0000000000001100", "1111111111101111", "0000000000011111", "0000000000011111", "0000000000000010", "0000000000000110", "0000000000100010", "1111111111110110", "1111111111011110", "0000000000000011", "0000000000010101", "0000000000011101", "1111111111100110", "1111111111011101", "1111111111101111", "1111111111101001", "1111111111111010", "1111111111101011", "1111111111001100", "0000000000000001", "1111111111110111", "1111111111010111", "1111111111101010", "0000000000001100", "0000000000100100", "1111111111101101", "1111111111010010", "0000000000011101", "0000000000100010", "0000000000000011", "1111111111100011", "0000000000000010", "0000000000011010", "0000000000001101", "0000000000010111", "1111111111101110", "0000000000010100", "0000000000100010", "1111111111110100", "0000000000001100", "1111111111110100", "1111111111000110", "1111111110111101", "1111111111100000", "0000000000000000", "1111111111100000", "1111111111010101", "0000000000000100", "1111111111110111", "0000000000000001", "1111111111011111", "0000000000010111", "0000000000011000", "0000000000010111", "0000000000000101", "1111111110111111", "1111111111010101", "1111111111010110", "0000000000001100", "0000000000001110", "0000000000010011", "1111111111011101", "1111111110101101", "1111111110110110", "0000000000010101", "1111111111100111", "1111111111001100", "1111111111100010", "0000000000100001", "0000000000011000", "1111111110110011", "1111111111101110", "0000000000001001", "0000000000011000", "0000000000011111", "1111111111000111", "1111111111011011", "1111111111110111", "1111111111111100", "0000000000000010", "1111111111001011", "1111111111011110", "0000000000001000", "1111111111100011", "0000000000000000", "1111111111010101", "1111111111100011", "0000000000101000", "1111111111010100", "0000000000110011", "1111111111111100", "0000000000100110", "0000000001010010", "0000000000001000", "0000000000010001", "1111111111001110", "0000000000111100", "0000000000000010", "1111111111110001", "0000000000001000", "1111111111011101", "1111111110111101", "1111111111100001", "1111111111110010", "1111111111101001", "1111111111110100", "0000000000101001", "0000000001000010", "0000000000010100", "0000000000011010", "0000000000011101", "0000000001010000", "0000000001000100", "0000000001001010", "1111111111011111", "0000000000110011", "0000000010010000", "0000000000110100", "0000000000000001", "1111111111101110", "0000000000001110", "1111111111001000", "1111111111010011", "0000000000101001", "1111111111100010", "1111111111010011", "1111111111001110", "1111111111001011", "1111111111110111", "0000000000010111", "1111111111001011", "1111111111100111", "1111111111111010", "0000000000000100", "1111111111101010", "1111111111101101", "1111111111011010", "1111111111100011", "1111111111010000", "1111111111101000", "0000000000001111", "1111111111101110", "1111111110111101", "1111111111101000", "0000000000111100", "0000000000011001", "0000000000000011", "1111111111111110", "0000000000100010", "0000000001000010", "0000000000010100", "0000000000000110", "1111111111110000", "0000000000111001", "0000000000010010", "0000000000110001", "0000000000101101", "1111111111100101", "1111111111100011", "1111111111001000", "1111111111001101", "0000000000000111", "1111111111101101", "1111111111001000", "1111111111101111", "1111111111100000", "1111111111101111", "1111111111100100", "0000000000100111", "0000000001000000", "0000000000001101", "1111111111110000", "0000000000001000", "0000000000110001", "1111111111111101", "0000000000000000", "1111111111010011", "0000000000100111", "1111111111111111", "1111111111001101", "0000000000111101", "0000000000000111", "1111111111110110", "1111111111111000", "1111111111110110", "1111111111011110", "1111111111110101", "0000000000001100", "0000000000000011", "1111111111111100", "1111111111111000", "1111111111110110", "1111111111110001", "0000000000011000", "1111111111110000", "0000000000000001", "1111111111010011", "1111111111111000", "1111111111110101", "1111111111001001", "1111111111110010", "1111111111111101", "1111111111111110", "1111111111010011", "0000000000000001", "0000000000111000", "0000000000010100", "0000000000000111", "0000000000001111", "1111111111101100", "1111111111011101", "0000000000010001", "1111111111100111", "0000000000001011", "1111111111111101", "1111111111011011", "0000000000000111", "1111111111110010", "1111111111101011", "1111111111111001", "0000000000000010", "1111111111001110", "1111111111011011", "1111111111101110", "1111111111111001", "1111111111010110", "0000000000000000", "1111111111100101", "0000000000000100", "0000000000001101", "0000000000101111", "0000000000000100", "1111111111111011", "0000000000001110", "0000000000001100", "1111111111011011", "1111111111110010", "1111111111011011", "1111111111011110", "1111111111010000", "1111111111101100", "1111111111011101", "1111111111001100", "1111111111011101", "1111111111000111", "1111111111111010", "1111111111010001", "1111111110110111", "1111111111011010", "0000000000011101", "0000000000001100", "1111111111001100", "1111111111000100", "0000000000000001", "0000000001000010", "1111111111010001", "0000000000000000", "0000000000000100", "1111111111110110", "1111111111110111", "0000000000000000", "1111111111110100", "1111111111001110", "1111111111101010", "0000000000101000", "0000000000011100", "1111111111111111", "1111111111011100", "0000000000001001", "0000000000111011", "0000000000000010", "1111111111111111", "0000000000010011", "0000000000001011", "1111111111101101", "0000000000001010", "0000000000000011", "0000000000001100", "1111111111101011", "1111111111111111", "0000000000010010", "1111111111001100", "0000000000000001", "1111111111111110", "0000000000011110", "1111111111100001", "1111111111010100", "0000000000001000", "1111111111101010", "0000000000001001", "0000000000001100", "0000000000000000", "1111111111101000", "1111111111010101", "0000000000100110", "0000000000100101", "0000000000010101", "0000000000010001", "1111111111000001", "0000000000000100", "0000000000010001", "0000000000100110", "0000000000101100", "0000000000001000", "0000000000011000", "1111111111000100", "1111111111010000", "1111111111010111", "0000000000001001", "1111111111110100", "1111111110111111", "1111111111011110", "1111111111110011", "1111111111100000", "1111111111001011", "1111111111111100", "1111111111011111", "1111111111100101", "1111111111101100", "1111111111101101", "1111111111110010", "0000000000001011", "1111111111110110", "0000000000110000", "0000000000110100", "1111111111101000", "1111111111010101", "1111111111100010", "0000000000011110", "0000000000001001", "0000000000000110", "1111111111100001", "1111111111001011", "1111111111110110", "0000000000000110", "1111111111001001", "1111111111011111", "0000000000000000", "0000000000000011", "0000000000001110", "1111111111001010", "1111111111100111", "1111111111101110", "1111111111101001", "0000000000000000", "1111111111000001", "1111111111010111", "0000000000011011", "0000000000001010", "0000000000000100", "1111111111010111", "1111111110111111", "0000000000010001", "0000000000110110", "0000000000110110", "1111111111100110", "1111111111101101", "1111111111110001", "0000000000010111", "0000000000011011", "1111111111100000", "1111111111100000", "1111111111100001", "1111111111011101", "0000000000001101", "1111111111110011", "1111111111011110", "1111111111100111", "1111111111111101", "1111111111110001", "0000000000001010", "0000000000000011", "0000000000000100", "0000000000001000", "0000000000010110", "1111111111111111", "0000000000110110", "0000000000110001", "1111111111101110", "0000000000100011", "1111111110100010", "1111111111011110", "0000000000000000", "0000000000000111", "1111111111111101", "1111111111100101", "0000000000001001", "0000000000001011", "1111111111101000", "0000000000000100", "0000000000011111", "1111111111110110", "0000000000011111", "0000000000010010", "0000000000000101", "0000000000000110", "1111111111011111", "0000000000011001", "0000000000001110", "1111111111011001", "0000000000001100", "1111111111111101", "1111111111100111", "0000000000001100", "0000000000101100", "1111111111110011", "1111111111111110", "1111111111010111", "0000000000001010", "0000000000000010", "0000000000010111", "1111111111110001", "1111111111110011", "1111111111101011", "0000000000000000", "0000000000111111", "0000000000001001", "0000000000000011", "0000000000010100", "1111111111100101", "0000000000000111", "1111111111101010", "0000000000001111", "0000000000011000", "0000000000000001", "1111111111100000", "1111111111111010", "0000000000000110", "0000000000000110", "1111111111111111", "0000000001111000", "0000000001101000", "0000000000100001", "0000000000000110", "0000000000001001", "0000000001100101", "0000000000001110", "0000000000011100", "1111111111110110", "1111111111110010", "0000000000101010", "0000000000001010", "0000000000011010", "1111111111100110", "1111111111011011", "1111111111011001", "1111111111111010", "1111111111100000", "1111111111001011", "1111111110111101", "1111111110110001", "1111111111001110", "0000000000000110", "1111111111101100", "1111111111101010", "1111111111010100", "1111111111000110", "1111111111011001", "0000000000000110", "0000000000000010", "1111111111110011", "0000000000000011", "0000000000110010", "0000000000001111", "0000000000000010", "1111111111000100", "1111111111100110", "0000000000100000", "0000000000001111", "0000000000001000", "1111111111011111", "1111111111100010", "0000000000000111", "0000000000010011", "1111111111111000", "0000000000000101", "1111111111010101", "0000000000001010", "0000000001001001", "0000000000110100", "0000000000001101", "0000000000010111", "0000000000010110", "1111111110111001", "1111111111111000", "0000000000011111", "0000000000000001", "1111111111101101", "1111111111101111", "1111111111100010", "0000000000010110", "1111111111110111", "1111111111111011", "0000000000000000", "0000000000000100", "1111111111000000", "0000000000010101", "0000000000001010", "1111111111100111", "0000000000000100", "1111111111100000", "0000000000001000", "1111111111100110", "1111111111111111", "1111111111011001", "0000000000100110", "0000000001000001", "1111111111010100", "0000000000100011", "0000000000111100", "0000000000000101", "0000000000011100", "1111111111111001", "0000000000000110", "0000000000011000", "1111111111010111", "1111111111101011", "0000000000010011", "1111111111110001", "1111111111100001", "1111111111101111", "1111111111101101", "1111111111100000", "1111111111110100", "1111111111010100", "1111111111110000", "1111111111010011", "0000000000111010", "0000000000100011", "1111111111000011", "1111111111101100", "1111111111000000", "0000000000010110", "0000000000111000", "0000000000111100", "1111111111100011", "0000000000000000", "0000000000110100", "0000000000110000", "0000000000000100", "1111111111111001", "1111111111111010", "1111111111101100", "1111111111101101", "1111111111101001", "1111111111101001", "1111111111101010", "1111111111011100", "1111111111010101", "0000000000000000", "0000000000011110", "1111111111100001", "1111111111010011", "1111111111000101", "1111111111101001", "0000000000010000", "1111111111101101", "0000000000001000", "1111111111111011", "1111111111100111", "1111111111101100", "1111111111100111", "1111111111110000", "1111111111111000", "0000000000001100", "0000000000000000", "1111111111100010", "1111111111111111", "0000000000100011", "1111111111111001", "1111111111110111", "1111111111101101", "0000000000011100", "0000000000001000", "0000000000000011", "1111111111111000", "1111111111010111", "1111111111111110", "1111111111111000", "0000000000000000", "1111111111100011", "1111111110111010", "1111111111010111", "1111111111011111", "1111111111010000", "1111111111100010", "1111111111010000", "1111111111110100", "0000000000001011", "0000000000011011", "1111111111100110", "1111111111111000", "0000000000001110", "0000000000110110", "0000000000101011", "1111111111110111", "1111111111100100", "1111111111010110", "1111111111101010", "1111111111010101", "1111111111101101", "0000000000000001", "1111111111010101", "1111111111111100", "1111111111110100", "0000000000001111", "1111111111010111", "1111111111000001", "1111111111110100", "1111111111011000", "1111111111100100", "1111111111001101", "1111111111011110", "0000000000000011", "0000000000110000", "1111111111110010", "1111111111101111", "0000000000001000", "0000000001000010", "0000000000001100", "0000000000000010", "0000000000000000", "1111111111101000", "1111111111011111", "1111111111001101", "0000000000000000", "1111111111101001", "1111111111001000", "1111111111010001", "1111111111111111", "0000000000010111", "1111111111100110", "1111111111000000", "1111111111011101", "1111111111000011", "1111111111110001", "1111111111101110", "1111111111110011", "0000000000000110", "1111111111101100", "0000000000010111", "0000000000000111", "0000000000010110", "1111111111111010", "0000000000001110", "1111111111111110", "0000000000010010", "1111111111110110", "1111111111110110", "0000000000000001", "0000000000011111", "1111111111100001", "1111111111100011", "1111111111110100", "0000000000000000", "1111111110011100", "1111111111010001", "0000000001010001", "0000000000111010", "0000000000100100", "1111111111000110", "0000000000001001", "0000000000101010", "0000000000010011", "1111111111100000", "0000000000010000", "0000000000000101", "1111111111110001", "1111111111111010", "1111111111110101", "0000000000000100", "1111111111110011", "1111111111101100", "1111111111011000", "1111111111100110", "1111111111111001", "1111111111001101", "1111111111010010", "1111111111010101", "1111111111101011", "0000000000000000", "0000000000101010", "0000000000011100", "0000000000001011", "0000000000011111", "1111111111101101", "0000000000010011", "0000000000001101", "1111111111111011", "0000000000101110", "0000000000001111", "1111111111101101", "1111111111101000", "1111111111000101", "0000000000011010", "1111111111110101", "0000000000000100", "1111111111111111", "1111111111011010", "0000000000010001", "1111111111110100", "1111111111011101", "1111111111101010", "1111111111101111", "0000000000000100", "0000000001010101", "0000000000100111", "0000000000011010", "0000000001000100", "0000000000001001", "1111111111110100", "0000000000011101", "0000000000100010", "0000000000000110", "1111111111001011", "1111111111111001", "0000000000000110", "0000000000000110", "1111111111100000", "1111111111110100", "1111111111101111", "1111111111101000", "1111111111011000", "0000000000100110", "0000000000011011", "1111111111100101", "1111111111111101", "1111111111110111", "0000000000010100", "0000000000001111", "0000000000000001", "1111111111010110", "1111111111001010", "1111111110101110", "1111111111111000", "1111111111010010", "0000000000101100", "1111111111100001", "1111111111001001", "0000000000010011", "1111111111010001", "1111111111111111", "1111111111111111", "0000000000001011", "0000000000011111", "0000000000000100", "1111111111011100", "1111111111111101", "0000000000110111", "1111111111110100", "0000000000001011", "0000000000001000", "0000000000010111", "1111111111110010", "0000000000011000", "0000000000000100", "1111111111101011", "0000000000011000", "0000000000010010", "0000000000110000", "0000000001011101", "0000000000101000", "0000000000100101", "0000000001001010", "0000000000011010", "0000000001010010", "0000000000010010", "0000000000000010", "0000000000101000", "1111111111110111", "0000000001001010", "1111111111110000", "1111111111110011", "1111111111111101", "1111111111101000", "0000000000111110", "1111111111010011", "1111111110100110", "1111111111001000", "1111111111001100", "0000000000101111", "0000000000010000", "1111111111100110", "1111111111010010", "1111111111111001", "0000000000011101", "1111111111011101", "1111111111011101", "1111111111011111", "0000000000000010", "1111111111011010", "1111111111001011", "1111111111101110", "1111111111100110", "1111111111101010", "1111111111110100", "1111111110111001", "1111111111110011", "0000000000000111", "0000000000011101", "1111111111100000", "1111111111001101", "1111111110110001", "0000000000000000", "0000000000010110", "0000000000100011", "0000000000000110", "1111111111111101", "1111111111101110", "1111111111100101", "0000000001011111", "1111111111111101", "1111111111011011", "1111111111100011", "1111111111101010", "0000000000101100", "1111111111111001", "1111111110111011", "1111111111101000", "1111111111100011", "0000000000011011", "1111111111011011", "1111111111011100", "0000000000010100", "0000000000001101", "1111111111110000", "1111111111101000", "1111111111101000", "1111111111010011", "0000000000001010", "1111111110111101", "1111111111101111", "1111111111110100", "1111111111001011", "1111111111110011", "1111111111100011", "0000000000000101", "1111111110111111", "1111111110110111", "0000000000001000", "1111111111010110", "0000000000000101", "1111111111100010", "1111111111011001", "0000000000001011", "1111111111101010", "0000000000011110", "1111111111001111", "0000000000101010", "0000000000100010", "1111111111101111", "1111111111110011", "1111111111111000", "0000000000011011", "0000000000111100", "0000000000000100", "0000000000011001", "1111111111011010", "1111111111011011", "1111111111000110", "1111111111011001", "0000000000100110", "1111111111101001", "1111111111100110", "1111111111100011", "1111111110100100", "1111111111100001", "1111111111001111", "1111111111111001", "1111111111101011", "1111111111010011", "1111111111111100", "1111111111111010", "0000000000110001", "0000000000011111", "1111111111101010", "1111111111110000", "1111111111100110", "1111111111111100", "0000000000011010", "0000000000000010", "0000000000110101", "0000000000000000", "1111111111011110", "1111111111011111", "0000000000010010", "0000000001110011", "0000000000100001", "1111111111111111", "1111111111011001", "0000000000000101", "0000000001001100", "0000000000100100", "1111111111011000", "0000000000011010", "1111111111100101", "0000000001101001", "0000000000011110", "1111111111110000", "0000000000000001", "1111111111010010", "0000000000001010", "0000000000101100", "0000000000011110", "1111111111111011", "1111111111100011", "1111111110010110", "1111111110100011", "1111111111100111", "0000000000000100", "1111111111001001", "1111111111011011", "1111111111101001", "1111111110101011", "0000000000111101", "0000000000000010", "0000000000100001", "1111111111100101", "0000000000000000", "0000000000100011", "0000000000110111", "0000000000001011", "1111111111001010", "0000000000001110", "0000000000010111", "0000000000101001", "1111111111011010", "1111111110111001", "1111111111111011", "1111111111000011", "0000000000000110", "0000000000011001", "0000000000100101", "1111111111100110", "1111111111010000", "0000000000100111", "0000000000011010", "0000000000001100", "1111111111110000", "1111111111111010", "1111111111001110", "1111111111101010", "1111111111100110", "0000000000101001", "0000000000100110", "1111111111100110", "1111111111011100", "0000000000010110", "1111111111110010", "1111111111101000", "1111111111110111", "1111111111101100", "1111111111111101", "1111111111101001", "1111111111001110", "0000000000011110", "1111111111100110", "1111111110101110", "1111111110100010", "1111111110101000", "1111111110110110", "1111111110010000", "1111111110000111", "1111111110101011", "1111111110010110", "1111111111111100", "1111111111001010", "1111111110110000", "1111111111000001", "1111111111101010", "0000000000001100", "0000000000011101", "1111111111111100", "1111111111110100", "1111111111100101", "0000000000010010", "0000000000000010", "0000000000100111", "1111111111111110", "0000000000110101", "1111111111110001", "1111111110110100", "1111111111011011", "0000000000010101", "1111111111100010", "1111111111001001", "1111111111101010", "0000000000010111", "0000000000000110", "1111111111011111", "1111111111101001", "1111111111100110", "1111111111111111", "1111111111101100", "0000000000001101", "0000000000111011", "0000000000001101", "0000000000101011", "0000000000101100", "1111111111111010", "0000000001010000", "1111111111101101", "1111111111111010", "0000000000000000", "1111111111111011", "1111111111100100", "1111111111111110", "1111111111110101", "1111111111101111", "1111111111110010", "1111111111011100", "0000000000001010", "1111111111011111", "0000000000011000", "1111111110101110", "0000000000010101", "1111111111110110", "1111111111101110", "1111111111010001", "1111111111100110", "0000000000010000", "1111111111011000", "0000000000101110", "0000000000111001", "1111111111110111", "0000000001001001", "1111111111111010", "1111111111111111", "0000000000011010", "1111111111111011", "1111111111101101", "0000000000110001", "0000000001000110", "0000000000111011", "0000000000100001", "0000000001100000", "0000000000110000", "0000000000001101", "0000000000000001", "1111111111010000", "0000000000000000", "1111111111110000", "1111111111111011", "1111111111100111", "1111111111101001", "1111111111010100", "1111111111111110", "0000000000000111", "1111111111110011", "1111111111010100", "1111111111011011", "1111111111111110", "0000000000001100", "0000000000000010", "1111111111001001", "1111111111011001", "1111111111000010", "1111111110110100", "1111111111100110", "1111111111101101", "1111111111010010", "1111111110111011", "1111111111011011", "0000000000011011", "0000000000110011", "1111111111001101", "1111111111001100", "0000000000101111", "0000000000101000", "0000000000011110", "1111111110100001", "1111111111101000", "0000000000000100", "1111111111110001", "1111111111100100", "1111111111111101", "0000000000011000", "0000000000011001", "0000000000001011", "1111111111010111", "0000000000011011", "1111111111010010", "1111111110111110", "1111111111110101", "0000000000011011", "1111111111101100", "1111111110111011", "0000000000011011", "1111111111111100", "1111111111010000", "0000000000100110", "0000000000111011", "1111111111101111", "1111111111111011", "1111111111111010", "0000000000011011", "0000000001001001", "0000000000100101", "1111111111100101", "1111111111111100", "0000000000010110", "0000000000101111", "0000000000010000", "0000000000100110", "1111111111000011", "0000000000001011", "0000000000010000", "0000000001100010", "0000000000111000", "1111111111111110", "0000000000011010", "0000000010001000", "0000000000110100", "1111111111101000", "1111111111101000", "1111111111000111", "1111111111010110", "1111111110110001", "0000000000010000", "1111111111110001", "1111111111010000", "1111111111000100", "1111111110110100", "1111111111111111", "1111111111010101", "0000000000010111", "0000000000001010", "1111111111001010", "1111111111110000", "1111111111000111", "0000000000100101", "0000000000000000", "1111111111011010", "1111111110110000", "0000000000011011", "1111111111111000", "1111111111011011", "1111111111000010", "0000000000000000", "0000000000110000", "1111111111110100", "1111111111001010", "1111111111111110", "0000000000100100", "0000000000010010", "1111111111010011", "0000000000100110", "0000000000101101", "0000000000101010", "1111111111101101", "1111111111100001", "0000000000000100", "0000000000001000", "0000000000010100", "1111111110111000", "0000000000001001", "0000000000100011", "1111111111011001", "0000000000001111", "1111111111001101", "1111111111111000", "1111111111110000", "0000000000010011", "0000000000100110", "1111111111101000", "1111111111011101", "0000000000000000", "0000000000011000", "0000000000100001", "1111111111010100", "1111111111101111", "1111111111011101", "1111111111111000", "0000000000000101", "1111111111001011", "0000000000000100", "0000000000010111", "1111111111111011", "1111111111010010", "1111111111110101", "1111111111011010", "1111111111011111", "1111111110101011", "1111111110101000", "1111111110111111", "1111111111110010", "1111111111010100", "1111111110111010", "1111111111010011", "1111111111101011", "1111111110111011", "1111111111100100", "1111111111000110", "1111111111110001", "1111111111010010", "0000000000001100", "0000000000010000", "1111111111110101", "1111111111011101", "1111111111011001", "0000000000110100", "0000000000101111", "0000000000011110", "0000000000010000", "0000000000100010", "1111111111110101", "1111111111111010", "1111111110100110", "1111111110101000", "1111111111011111", "1111111111011010", "1111111111100101", "1111111110111110", "1111111111000001", "1111111111001110", "1111111110110101", "1111111111000000", "1111111110110111", "1111111111101000", "0000000000000000", "1111111111001000", "1111111111101010", "1111111111111100", "1111111111100100", "1111111111001100", "1111111111111110", "0000000001010110", "0000000000111110", "0000000000011110", "1111111111100001", "0000000000010101", "0000000000001111", "1111111111010001", "1111111111010101", "1111111111011110", "0000000001001100", "0000000000110010", "1111111110111111", "1111111111000110", "1111111111100100", "0000000000011001", "1111111110111111", "1111111111010011", "0000000000010100", "0000000000000111", "0000000000100001", "1111111111100011", "0000000000000010", "0000000000001100", "0000000000000110", "0000000000000110", "0000000000011000", "0000000000111001", "0000000000100101", "0000000000010010", "1111111111111000", "0000000000000100", "1111111111010100", "1111111111111110", "0000000000101100", "1111111111001101", "1111111111001001", "1111111111111000", "0000000000010001", "0000000000100100", "1111111110111111", "1111111111110111", "0000000000001110", "1111111111101101", "1111111111001110", "1111111111101000", "0000000000000001", "0000000000001111", "1111111110111010", "1111111111001111", "1111111111110111", "0000000000010011", "0000000000000100", "1111111111110110", "1111111111110010", "0000000000000001", "0000000000100000", "1111111111111011", "1111111111100111", "1111111111000100", "0000000001010000", "1111111111110110", "0000000000010011", "1111111111010010", "0000000000100110", "0000000001011000", "0000000000011011", "1111111111101101", "1111111111000001", "0000000000100001", "0000000000110111", "1111111111100001", "1111111111010010", "0000000000000011", "0000000000100101", "0000000001000010", "1111111111011111", "1111111111100000", "0000000000001100", "1111111111100011", "0000000000100001", "0000000000001011", "0000000000111110", "1111111111111110", "0000000000001001", "0000000000010011", "0000000000111001", "1111111111100110", "0000000000101000", "0000000000100100", "0000000000011011", "1111111111010110", "0000000000001000", "0000000001001101", "0000000000000011", "1111111111000100", "1111111111100110", "1111111111101010", "0000000000010110", "0000000000001100", "1111111111100100", "1111111111111011", "1111111111111110", "0000000000010111", "0000000000000110", "1111111111110101", "0000000000000010", "0000000000010110", "1111111111111011", "1111111110101101", "0000000000001010", "0000000000001100", "0000000000100110", "1111111111010111", "1111111111010011", "0000000001101011", "0000000001000001", "0000000000000100", "1111111110101000", "1111111111011000", "1111111111111011", "1111111111010111", "1111111111011011", "1111111110110010", "0000000000000111", "1111111111001001", "1111111111001111", "1111111110111111", "1111111111010011", "1111111111010100", "1111111111111111", "0000000000010101", "0000000001101010", "1111111111010110", "1111111111101010", "1111111111111111", "0000000001011101", "0000000000001001", "1111111111010110", "0000000000100010", "1111111111011000", "1111111111111011", "1111111111011110", "1111111111111110", "0000000001010110", "1111111111110010", "1111111110111100", "1111111111100001", "0000000000011100", "0000000000111111", "1111111111010100", "1111111110101101", "1111111111010001", "0000000000010110", "0000000000011000", "0000000000000110", "1111111111110011", "1111111111011011", "0000000000001110", "0000000000100001", "0000000000001001", "0000000000010101", "1111111111010101", "1111111111011111", "1111111111110011", "0000000000110100", "1111111111110111", "0000000000010011", "0000000000001001", "1111111111001111", "0000000000100010", "0000000000001010", "0000000000000000", "1111111111111100", "1111111111101001", "0000000000100101", "0000000000000000", "1111111111111111", "0000000000000101", "0000000000010001", "0000000000001001", "1111111111101101", "0000000000001100", "1111111111101100", "0000000000100011", "0000000000000000", "0000000000010010", "1111111111100101", "1111111111101111", "0000000000000111", "1111111111110110", "0000000000000000", "1111111111101001", "1111111111100100", "0000000000000100", "0000000000110001", "0000000000010000", "1111111111100011", "1111111111011110", "0000000000000111", "0000000000111100", "1111111111101000", "1111111111010100", "1111111111110001", "0000000000011000", "1111111110111110", "1111111110000011", "1111111111101101", "1111111111100100", "1111111111001011", "1111111111000011", "1111111111101011", "0000000000000111", "1111111111100001", "1111111111000111", "1111111111010100", "0000000000100110", "0000000000101001", "0000000000000000", "1111111110011011", "0000000001001100", "0000000000110101", "1111111111011111", "1111111111001011", "1111111111111010", "0000000000010000", "1111111111110100", "1111111111011100", "1111111111001001", "0000000000001110", "0000000000101001", "0000000000000011", "1111111111011101", "1111111110110100", "1111111111001100", "1111111111110001", "1111111111011111", "1111111111010110", "1111111111010000", "1111111111100011", "0000000001110000", "0000000000011000", "1111111111110000", "1111111111100101", "1111111111011010", "0000000000100001", "1111111111100000", "1111111111110000", "1111111111010110", "1111111111001110", "0000000000110111", "1111111111111100", "1111111111101100", "0000000000000000", "1111111111001100", "0000000000011011", "1111111111010100", "1111111111100001", "0000000000000100", "0000000000000011", "0000000000000101", "1111111111011111", "0000000000100011", "0000000000011101", "1111111111010001", "0000000000011001", "1111111111011110", "1111111111111101", "1111111111101101", "1111111111011111", "1111111111101001", "1111111111110000", "1111111111001011", "1111111110110100", "1111111111101000", "1111111110110101", "1111111111000010", "1111111111001110", "1111111111100011", "0000000000000110", "1111111110100011", "1111111110011001", "1111111111111110", "0000000000000011", "1111111111010011", "0000000000010001", "1111111111111101", "0000000000110001", "1111111111100111", "1111111111100111", "0000000001001010", "0000000001001001", "0000000000000101", "1111111111101101", "1111111111101011", "0000000000010111", "0000000000100000", "1111111111011101", "0000000000000011", "0000000000001100", "1111111111011001", "1111111111001001", "1111111111110001", "0000000000001011", "0000000000010011", "1111111111101101", "1111111111101111", "1111111111000101", "1111111111010111", "1111111111101000", "0000000000110011", "0000000000011001", "1111111111111101", "1111111111110000", "0000000000101111", "0000000000110011", "0000000000010100", "0000000000001111", "0000000000001010", "1111111111110011", "0000000000001100", "0000000000001101", "0000000000010110", "0000000000010011", "0000000000100001", "0000000000011111", "1111111111111011", "1111111111101000", "1111111111111110", "0000000000010011", "1111111111111101", "0000000000100101", "0000000000000000", "0000000000011101", "1111111111011000", "1111111111001001", "1111111111110011", "1111111111101110", "1111111111111000", "1111111111100111", "0000000000011111", "1111111111101111", "1111111111011100", "1111111111100010", "0000000000101010", "0000000000101000", "0000000000001100", "1111111111011100", "0000000000010001", "0000000000100001", "0000000000000100", "1111111111111110", "0000000000110101", "0000000000011111", "1111111111011001", "1111111111110110", "1111111111111100", "0000000000001001", "0000000000010010", "1111111111101111", "0000000000011011", "0000000000001011", "0000000000000000", "0000000000010111", "0000000000011000", "0000000001010101", "1111111111100100", "1111111110111110", "1111111111100011", "0000000000010010", "0000000000011111", "1111111111001001", "1111111110100001", "1111111111010110", "1111111111111111", "1111111111101111", "1111111111101100", "1111111110101001", "1111111111010110", "0000000000011011", "0000000000000001", "0000000000001010", "1111111111111110", "1111111111111010", "1111111111111010", "0000000000001000", "0000000000000011", "1111111111011000", "0000000000010000", "0000000000100111", "0000000000101011", "1111111111111100", "1111111111000110", "1111111111111110", "0000000000000111", "0000000000110111", "0000000000100010", "1111111110100110", "1111111111001110", "0000000000010100", "0000000000011100", "0000000000101000", "1111111111110110", "1111111110111011", "1111111111100000", "1111111111010110", "1111111111011001", "1111111111111100", "1111111111001000", "0000000000000011", "1111111110100001", "1111111111010010", "1111111110111011", "1111111111111010", "1111111111110000", "1111111111010010", "1111111111111111", "1111111111101000", "1111111111111001", "1111111111100111", "1111111111110010", "1111111111100001", "0000000000010111", "1111111111100111", "1111111111110101", "0000000000000111", "1111111111011010", "0000000000001111", "0000000000000010", "0000000001001111", "0000000000101010", "0000000000001011", "1111111111000000", "1111111111011001", "1111111111110010", "0000000000110100", "1111111111010100", "1111111111011010", "0000000000001101", "0000000000100010", "0000000000101010", "1111111111101011", "1111111111111011", "0000000000010001", "0000000000000111", "1111111111100000", "1111111111101111", "1111111111000000", "1111111111001000", "1111111111011111", "1111111111001001", "1111111111001110", "1111111110010111", "1111111111001001", "1111111111001100", "1111111111111000", "0000000000000111", "0000000001000111", "0000000000000000", "1111111111111111", "0000000000001010", "0000000000111001", "0000000000001110", "0000000000000010", "0000000000001111", "1111111111011101", "0000000001010001", "0000000000111000", "1111111111101010", "0000000000000010", "1111111111101001", "1111111111111100", "0000000000110000", "0000000000101001", "0000000000011100", "1111111111100011", "1111111111100101", "0000000000010111", "0000000001001011", "0000000000011011", "1111111110101101", "1111111111101010", "1111111111010011", "1111111111011001", "1111111111110101", "1111111110101101", "1111111111000111", "1111111111001101", "1111111111001100", "1111111111110101", "1111111111001010", "1111111110001110", "1111111110101110", "0000000000010001", "1111111111100001", "0000000000000100", "1111111111101110", "1111111111100110", "0000000000011000", "1111111111110000", "0000000001101001", "0000000001001011", "0000000000011101", "0000000001010001", "0000000001000011", "1111111111100000", "1111111111110110", "0000000000101000", "0000000001010011", "0000000000010011", "1111111111100000", "0000000000010101", "0000000000001110", "1111111111101111", "1111111111010110", "1111111111101001", "1111111111110001", "1111111111100000", "1111111111101001", "1111111111100010", "1111111111001001", "1111111111011110", "1111111111111100", "0000000000011011", "0000000000101110", "1111111111010101", "1111111111011110", "1111111111111100", "0000000000001011", "0000000000110000", "1111111111111001", "1111111111100111", "1111111111100101", "1111111111100110", "1111111111000111", "0000000000010101", "0000000000001011", "1111111111000101", "1111111111100100", "0000000000000011", "0000000000000110", "0000000000010000", "0000000000001001", "1111111111100110", "0000000000011100", "0000000000000101", "0000000000001101", "0000000000000001", "1111111111011010", "1111111111100000", "1111111111101011", "1111111111101001", "0000000000001001", "1111111111111000", "1111111111100101", "1111111111101110", "1111111111011000", "1111111111101001", "0000000000001001", "0000000000000011", "1111111111001100", "1111111110111101", "1111111111101000", "0000000000101001", "0000000000011000", "1111111111100000", "0000000000000001", "1111111111101000", "1111111111101000", "1111111111111100", "1111111111110001", "0000000000111001", "0000000000010010", "0000000000110010", "0000000000001011", "0000000000111110", "0000000000101001", "0000000000101110", "0000000000011001", "1111111111111000", "1111111111000101", "1111111110111101", "1111111111001001", "1111111111111100", "1111111111110111", "1111111111110000", "1111111111110011", "1111111111111111", "0000000000011100", "0000000000001001", "1111111111101111", "0000000000010101", "1111111111110001", "0000000000001001", "1111111111110110", "1111111111101011", "1111111111111000", "0000000000000111", "0000000000010001", "1111111111111111", "0000000000011000", "0000000000011101", "0000000000111110", "0000000001001011", "0000000000000110", "1111111111101111", "1111111110111100", "1111111111100101", "1111111111000100", "1111111111011111", "1111111111101000", "0000000000000000", "1111111111110001", "0000000000000110", "1111111111111010", "1111111111001110", "0000000000011111", "1111111111111010", "1111111111111101", "1111111111011110", "1111111111011010", "1111111111100110", "0000000000000100", "0000000000000100", "1111111111011000", "1111111111101111", "1111111111011010", "1111111111101101", "1111111111101100", "1111111111101001", "1111111111101001", "0000000000001101", "0000000001010100", "0000000001101010", "0000000001000100", "0000000000000000", "0000000000000010", "0000000000010010", "0000000000001100", "1111111111101110", "1111111111101111", "1111111111011100", "1111111110110110", "1111111111100011", "1111111111110000", "1111111111111110", "1111111111101010", "1111111111011000", "1111111111010110", "1111111111110101", "0000000000101001", "0000000000101010", "0000000000010010", "1111111111110011", "1111111111101110", "1111111110110101", "1111111111001000", "1111111111011010", "0000000000100010", "0000000000110001", "1111111111000101", "1111111111001101", "1111111110111101", "1111111111011011", "1111111111110110", "0000000000000111", "0000000000000011", "1111111111111111", "1111111111100101", "0000000000100101", "0000000001000101", "0000000000101110", "0000000000011000", "1111111111110011", "0000000000000011", "1111111111110100", "1111111111001111", "1111111111101111", "1111111111011101", "1111111111111111", "1111111111110001", "0000000000000001", "0000000000011010", "1111111111111100", "1111111111010011", "0000000000000100", "0000000000011110", "0000000001100001", "1111111111111001", "1111111111101101", "1111111111110101", "0000000001000001", "0000000000001110", "0000000000110110", "0000000000101011", "1111111111100010", "0000000000010101", "0000000000011100", "0000000000111010", "0000000000101100", "1111111111010001", "1111111111111110", "1111111111110000", "1111111111100001", "1111111111110111", "1111111111010011", "1111111111100001", "0000000000001001", "1111111111101010", "0000000000011000", "1111111111011001", "1111111111101110", "0000000000101100", "0000000000101011", "1111111111110010", "1111111111110011", "1111111111110111", "0000000000100110", "1111111111100100", "1111111111001011", "0000000000001110", "0000000000110001", "0000000000000000", "0000000000010011", "1111111111100101", "0000000000001111", "0000000000011010", "0000000000110100", "1111111111111001", "0000000000000001", "1111111111101100", "1111111111100101", "0000000000000111", "1111111111111010", "1111111111110000", "0000000000000001", "0000000001000001", "0000000000110000", "1111111111101100", "1111111111011010", "0000000000110001", "0000000001101000", "0000000000010001", "1111111111111100", "1111111111110111", "1111111111111011", "0000000001010000", "0000000000000110", "1111111111101100", "1111111111010001", "1111111111100110", "0000000000101001", "1111111111110100", "1111111111010101", "1111111111001010", "1111111111111100", "1111111111101001", "1111111111111010", "1111111111110001", "1111111111001011", "1111111111110101", "1111111111000110", "1111111111010001", "1111111111010110", "1111111110111000", "0000000000001001", "1111111111110101", "1111111111011100", "1111111111110111", "1111111111010000", "0000000000000001", "0000000000010101", "1111111111010001", "1111111111000100", "1111111111011000", "0000000000101001", "0000000000000110", "1111111111101011", "1111111111000111", "1111111111011101", "1111111111001100", "1111111111111000", "1111111111101111", "1111111111100000", "1111111111100111", "1111111111101001", "1111111111100110", "1111111111100110", "1111111111101000", "1111111111000110", "1111111111100000", "0000000000011100", "1111111111010101", "1111111111110010", "1111111111100111", "1111111111011001", "0000000000101010", "0000000000011011", "1111111110111010", "1111111110111010", "0000000000011000", "0000000000000000", "0000000000011001", "1111111111110001", "1111111111100011", "1111111111001110", "1111111111100100", "1111111111101010", "1111111111001010", "1111111111001111", "1111111111100001", "1111111111100100", "1111111111000011", "1111111111101000", "1111111111110111", "1111111111010000", "1111111111110101", "1111111111111100", "0000000000100101", "0000000000001101", "1111111110011100", "1111111111001101", "0000000000000100", "0000000000010000", "1111111111111011", "1111111111101001", "1111111111101100", "0000000000100010", "0000000000110010", "0000000000010010", "0000000000010010", "0000000000010101", "0000000000000101", "0000000000000100", "0000000000001010", "1111111111101110", "0000000000010111", "0000000000001110", "0000000000001110", "0000000000001000", "1111111111010010", "1111111111111110", "1111111111111010", "1111111111101000", "1111111111001111", "0000000000001011", "1111111111011011", "1111111111110110", "1111111111110110", "0000000000001000", "0000000000011010", "1111111111110000", "0000000000001111", "1111111111011011", "1111111111101011", "1111111110101001", "1111111111101001", "1111111111110100", "1111111111010110", "1111111111100011", "1111111111011001", "1111111110110111", "0000000000000110", "0000000000000100", "1111111111011010", "1111111111101100", "1111111111001011", "0000000001001010", "0000000000010000", "0000000000000011", "0000000001000100", "1111111111101001", "0000000000001010", "0000000001000010", "0000000000011000", "0000000000000000", "1111111111110100", "0000000000011111", "0000000000011111", "0000000000010001", "1111111111000110", "0000000000000100", "1111111111000111", "1111111110101100", "1111111111010110", "1111111111111011", "1111111111110111", "0000000000100111", "1111111111100000", "1111111111111110", "1111111111110010", "0000000000001110", "0000000000010100", "1111111111011000", "1111111111110011", "1111111111011110", "1111111111100111", "0000000000010110", "1111111111001011", "1111111111111110", "1111111111010111", "1111111111110010", "1111111111100110", "0000000000001101", "0000000001010110", "1111111111111100", "0000000000000001", "1111111111000110", "1111111111000111", "0000000000010110", "0000000000000110", "1111111111110101", "1111111111100110", "1111111111000001", "1111111110010110", "0000000000110100", "0000000001011000", "0000000001000100", "0000000000001101", "1111111111110000", "0000000000111100", "1111111111110100", "0000000000000001", "0000000000001100", "1111111111111011", "1111111111001011", "1111111111001100", "1111111111001100", "1111111111111000", "0000000000010000", "0000000000000010", "0000000000000000", "0000000000000101", "0000000000111001", "1111111111010001", "1111111110111101", "1111111110111011", "1111111111001110", "1111111111101110", "1111111111001001", "1111111110111000", "1111111110111011", "1111111111010111", "1111111111001000", "1111111111011101", "1111111110110011", "1111111111110000", "0000000000000001", "1111111111101101", "1111111111110000", "0000000000011110", "0000000000111001", "1111111111111101", "1111111111110001", "1111111111101111", "0000000001001101", "0000000000010001", "0000000000110110", "0000000000001010", "1111111111011101", "1111111111000100", "1111111111110110", "0000000000011000", "0000000000111010", "0000000000011000", "1111111110111011", "1111111111001111", "1111111111100000", "0000000000000101", "0000000000010000", "1111111111110011", "1111111111110100", "1111111111110111", "1111111111010111", "1111111111110101", "1111111111101010", "0000000000010111", "1111111111010000", "0000000000000000", "1111111111111111", "0000000000011010", "0000000000110100", "0000000000001100", "0000000000011101", "0000000000010100", "1111111110011010", "1111111111011001", "1111111111100111", "0000000000011010", "0000000000100011", "1111111111010010", "1111111110100010", "1111111111000010", "1111111111010110", "0000000000001001", "0000000000000011", "1111111111101011", "1111111111100000", "1111111111110000", "1111111111101011", "1111111111110101", "0000000000010011", "1111111111101101", "0000000000000101", "0000000000010110", "0000000000101100", "0000000000101101", "0000000000001111", "0000000000001011", "0000000001000011", "1111111111000000", "1111111111011101", "1111111111110010", "0000000000011000", "0000000001000001", "1111111111101111", "1111111111011111", "1111111110011100", "1111111110110111", "1111111111001000", "0000000000110011", "0000000000001100", "1111111111101110", "1111111111001111", "1111111110110101", "0000000000100111", "0000000000010101", "0000000000011011", "0000000000000101", "0000000000010100", "1111111111101110", "1111111111011110", "1111111111100011", "1111111111110000", "0000000000011010", "1111111111100011", "0000000000011011", "1111111111111011", "1111111111110011", "1111111111111010", "0000000000110111", "0000000000101100", "0000000000011110", "0000000000101000", "0000000001001101", "0000000001011100", "1111111111100001", "1111111111011010", "0000000000001000", "0000000000011110", "1111111111101100", "1111111111111001", "1111111111010001", "1111111111111101", "0000000000010111", "1111111111010000", "1111111111111010", "1111111111110010", "1111111111101110", "0000000000000100", "0000000000010010", "1111111111001110", "1111111111101110", "1111111110111110", "1111111110101110", "0000000000101010", "0000000000001001", "0000000001001010", "0000000000010000", "1111111110111100", "1111111111110110", "0000000000001111", "0000000000101011", "0000000000110010", "1111111111001001", "1111111111010101", "1111111111000100", "0000000000111000", "0000000001010000", "1111111111010101", "0000000000110101", "0000000000000111", "1111111111111100", "1111111111000100", "0000000000010000", "1111111111101001", "1111111111100010", "1111111111010101", "1111111111000110", "1111111111110001", "1111111111111000", "0000000000000011", "1111111111011100", "1111111110110001", "1111111101111110", "0000000000011011", "1111111111001000", "1111111111101100", "1111111111110001", "1111111111010011", "1111111111111101", "1111111111111110", "0000000000011000", "1111111111111010", "1111111111011000", "1111111110111011", "1111111111001111", "1111111111100101", "1111111111101001", "1111111111011010", "0000000000001010", "0000000000110101", "0000000000110011", "0000000001000101", "0000000000010110", "0000000000100000", "1111111111110110", "0000000000011001", "0000000000011100", "1111111111101101", "0000000000000000", "1111111111100101", "1111111110111010", "1111111111000011", "1111111111011110", "0000000000000001", "1111111111010001", "1111111111101010", "0000000000000110", "1111111111101011", "1111111111110011", "1111111111010110", "1111111111010000", "1111111111110101", "0000000000001100", "1111111111101010", "0000000000010010", "0000000000011100", "1111111111011100", "1111111111111110", "0000000000100011", "0000000000111110", "0000000000000010", "1111111111101111", "1111111111110000", "1111111111110110", "1111111111110100", "0000000000110111", "0000000000100010", "1111111111110100", "1111111111111111", "1111111111111001", "0000000000011010", "1111111111000011", "1111111111010100", "1111111111101001", "1111111110111110", "1111111111101101", "0000000000001010", "1111111111110111", "1111111111000110", "1111111111110100", "1111111111110110", "0000000000001100", "0000000000010010", "0000000000110001", "1111111111111011", "0000000000111010", "0000000000010111", "0000000000101000", "0000000000001011", "1111111111111001", "0000000000111010", "0000000000011110", "0000000000011001", "1111111111011010", "1111111111100010", "1111111111011111", "1111111111101010", "1111111111001011", "1111111111110001", "1111111111000111", "1111111111010010", "1111111111101111", "1111111111100110", "1111111111001111", "1111111111011010", "1111111111001001", "1111111111010001", "0000000000000110", "0000000000100000", "0000000000011011", "0000000000110100", "0000000000001000", "0000000000100110", "1111111111111001", "1111111111011000", "0000000001010101", "0000000000111011", "0000000000011001", "1111111111101001", "1111111111010111", "1111111111010111", "1111111111101001", "0000000000000010", "0000000000001010", "1111111111100010", "1111111111100100", "1111111110110001", "1111111111001110", "1111111111010011", "1111111111101010", "1111111111001110", "1111111111111110", "1111111111000110", "0000000000111101", "0000000000110111", "1111111111111010", "1111111111100000", "1111111111101111", "0000000000111100", "0000000000011101", "1111111111011101", "0000000000000001", "0000000000000110", "1111111111101100", "1111111111011000", "1111111111101110", "0000000000000111", "0000000000100010", "1111111111011010", "1111111111111000", "1111111111101101", "1111111111111100", "0000000000100000", "1111111111111110", "0000000000100010", "0000000000100101", "0000000000010110", "1111111111110010", "0000000001000110", "0000000000101010", "0000000000010000", "0000000000110101", "1111111111111111", "0000000000000001", "0000000000000000", "1111111111011000", "1111111111010101", "1111111111100110", "0000000000011000", "1111111111110010", "1111111111010001", "1111111111000000", "1111111111001000", "1111111111101011", "1111111111111000", "1111111111111101", "1111111111011001", "0000000000000101", "1111111111010010", "1111111111010101", "1111111111111110", "0000000000111010", "0000000000000101", "0000000000000001", "1111111111101001", "1111111111110111", "0000000000100011", "0000000000001001", "1111111111100110", "1111111111110001", "1111111110111100", "1111111111110000", "1111111111101011", "1111111111011100", "1111111111111000", "1111111110010111", "1111111110110001", "1111111110100010", "0000000000000000", "1111111111100111", "1111111111011111", "1111111111001101", "1111111111101011", "0000000000110111", "0000000000010111", "1111111111110101", "1111111111001111", "1111111111011100", "0000000000110100", "0000000000100110", "1111111111101101", "1111111110011100", "0000000000001011", "0000000001000000", "0000000000100011", "1111111111111000", "1111111111111101", "1111111111110110", "1111111111011000", "1111111111111110", "1111111111111100", "0000000000110110", "0000000000010011", "1111111111010100", "1111111111011011", "1111111111100001", "0000000000010011", "0000000000100010", "1111111110111100", "1111111111000110", "1111111111100000", "0000000000000111", "1111111111100110", "0000000000000111", "0000000000000101", "1111111111011101", "1111111111011001", "0000000000001111", "0000000000010110", "0000000000001101", "1111111111110010", "1111111111101101", "1111111111110010", "0000000000011001", "1111111111111010", "0000000000001101", "0000000000100100", "1111111111000001", "1111111111101001", "0000000000110100", "0000000000111010", "1111111111100101", "1111111111101000", "0000000000000011", "0000000000001111", "0000000000111110", "0000000000010000", "0000000000000101", "1111111111010111", "0000000000001011", "0000000000001101", "0000000000000000", "1111111111101011", "1111111111011010", "1111111110111011", "1111111111100111", "0000000000110001", "0000000000011001", "1111111111000001", "1111111111110110", "1111111110110110", "1111111111010101", "0000000000001101", "1111111111111001", "1111111111001010", "1111111110111100", "1111111111011110", "1111111111110011", "0000000000011101", "0000000000001011", "1111111111110111", "1111111110110001", "1111111110010101", "0000000000010000", "0000000000011010", "0000000001000001", "1111111111101101", "1111111111011010", "1111111111001001", "1111111111100001", "0000000001000100", "0000000001110011", "0000000000101010", "1111111111010111", "1111111111000111", "1111111110101010", "0000000000000101", "0000000000100100", "0000000000000011", "0000000000001001", "1111111111101000", "1111111111010111", "1111111111100010", "1111111111111100", "0000000000000110", "0000000000001101", "1111111111110111", "1111111110010100", "1111111111011100", "1111111111011100", "0000000000011111", "0000000000001000", "1111111111101010", "1111111111001001", "1111111111000111", "0000000000001111", "0000000001001100", "0000000000010111", "1111111111100110", "1111111110110001", "1111111111011101", "1111111111110000", "0000000000101100", "0000000000001110", "1111111111101111", "0000000000101011", "0000000000011110", "1111111111111110", "1111111111100000", "1111111110110011", "1111111111111000", "0000000000010001", "0000000000000100", "1111111111001011", "1111111110111000", "1111111110111111", "0000000000000110", "0000000000010011", "1111111111110010", "1111111111101010", "0000000000011010", "0000000000000000", "0000000000001100", "0000000000000111", "1111111111111011", "1111111111111010", "1111111111110100", "0000000000011010", "1111111111000111", "1111111111010001", "1111111111100101", "0000000000010110", "0000000000000111", "1111111111111000", "1111111111011110", "1111111110101011", "1111111111100110", "1111111110111110", "0000000000010000", "1111111111101010", "1111111111001001", "1111111111001000", "1111111111010000", "1111111111101011", "1111111111110001", "1111111111011100", "1111111111001011", "1111111111100001", "1111111111011110", "0000000000011101", "0000000000010100", "1111111111011110", "1111111111011001", "0000000000001110", "0000000000001101", "0000000000011010", "0000000000011101", "1111111111011101", "0000000000000111", "1111111111011011", "0000000000101110", "0000000000101111", "1111111111110000", "1111111111110110", "1111111111011110", "1111111111111100", "0000000000111100", "0000000000101011", "1111111111110100", "0000000000000101", "1111111111110000", "1111111111000110", "0000000000000010", "0000000000010110", "0000000000010100", "1111111110111110", "1111111110111011", "1111111110010100", "1111111111100000", "1111111111110011", "0000000000110001", "0000000001000000", "0000000000000000", "1111111111100010", "1111111111010010", "0000000000010101", "0000000000000000", "0000000000010001", "1111111111100100", "1111111111011010", "1111111111110000", "1111111111111101", "0000000000001010", "0000000000010001", "1111111111111100", "1111111110111011", "1111111111010101", "0000000000010101", "0000000000011011", "1111111111100000", "1111111111111111", "1111111111101001", "1111111111110100");
    Plus112_i_1 <= ("1111111111110111", "1111111111010011", "1111111110010110", "1111111111111111", "0000000000000011", "1111111111101101", "1111111110111110", "1111111110111100", "1111111111001110", "1111111111011110", "1111111111001001", "1111111111010011", "1111111111001100", "1111111111011100", "1111111111100101", "1111111111101011");
    Times212_i_1 <= ("0000000000011111", "1111111111110111", "0000000000111100", "1111111111001000", "0000000001000101", "1111111110111011", "0000000000110101", "1111111111011101", "1111111111100010", "0000000000100000", "0000000010000100", "1111111110100001", "0000000000001111", "1111111110001010", "0000000000011100", "0000000001011101", "0000000000000001", "1111111111001101", "0000000000011001", "1111111111100111", "1111111111100100", "1111111111010001", "0000000000000000", "1111111111110000", "0000000000101001", "0000000000010001", "1111111111001011", "1111111111011001", "0000000001110011", "1111111111010011", "1111111111111110", "0000000000000001", "0000000000000001", "0000000000000010", "0000000000010111", "1111111111101010", "0000000000001111", "1111111111011100", "1111111111100001", "1111111111111001", "1111111110111111", "1111111111111111", "0000000001100110", "1111111110100111", "0000000000100111", "1111111111111010", "1111111110011010", "0000000001011001", "1111111111011111", "0000000001001100", "1111111110111110", "0000000001000001", "1111111111110111", "0000000000001010", "0000000000110100", "1111111110101101", "1111111111001001", "0000000000010110", "0000000001011110", "1111111111110000", "0000000000001000", "1111111111111000", "0000000010000100", "0000000000001010", "1111111111010000", "1111111111111010", "1111111110111110", "1111111110101100", "1111111111001000", "0000000001100101", "0000000000011010", "1111111111011111", "0000000000100001", "0000000000000100", "0000000000010001", "1111111111110110", "1111111111100111", "1111111111111000", "1111111111111010", "0000000000001110", "1111111111100101", "0000000000010100", "0000000001000101", "1111111111100010", "1111111110100000", "0000000001101111", "0000000000010000", "1111111111010000", "0000000001000011", "1111111110110110", "0000000000000011", "1111111110100001", "0000000000001000", "0000000001000111", "0000000000100001", "1111111111110111", "1111111101111110", "0000000000000001", "0000000000010001", "0000000001000010", "0000000000110111", "0000000000001110", "0000000000000101", "0000000001100101", "1111111111010001", "0000000001000100", "1111111111101111", "1111111110110001", "1111111111001111", "1111111111010101", "0000000000011011", "0000000000100010", "1111111111100100", "1111111111110001", "1111111111101111", "1111111111110010", "1111111111100111", "1111111111111101", "1111111111101110", "0000000000001001", "0000000000010001", "1111111111110001", "1111111111111000", "0000000000000000", "0000000000000101", "0000000000010001", "0000000000001101", "1111111111010100", "0000000000001100", "1111111111101000", "1111111111011101", "1111111111100010", "1111111111111111", "0000000001100100", "1111111111000000", "0000000000001101", "0000000000011011", "1111111111000100", "0000000000100101", "1111111111011011", "1111111111001111", "1111111111111100", "0000000000101011", "0000000001000001", "1111111111010100", "0000000000101101", "1111111111100010", "0000000000011101", "0000000000001010", "1111111111100110", "1111111111011100", "0000000000001111", "1111111111100000", "1111111111100011", "1111111111110011", "0000000000000001", "1111111111110110", "1111111111101110", "1111111111111011", "0000000000011001", "1111111111010111", "0000000001110111", "1111111111010010", "1111111111100111", "0000000000000101", "1111111111111110", "0000000000000111", "0000000000110000", "0000000000000000", "1111111111001101", "0000000000100011", "1111111111101001", "0000000000011111", "1111111110110111", "0000000000010011", "1111111111010101", "0000000000100001", "1111111111011010", "0000000000101100", "1111111111011111", "1111111111111001", "0000000001000100", "0000000000001111", "1111111111010001", "1111111111010111", "0000000000100100", "1111111111110101", "0000000000001110", "1111111111101111", "0000000000101001", "0000000000000100", "1111111111100010", "1111111111101000", "1111111111010110", "0000000000101110", "0000000000100111", "1111111111101110", "1111111111101011", "1111111111110010", "1111111111101000", "1111111111011000", "0000000001100111", "1111111110101010", "0000000000111011", "0000000001111001", "1111111110001111", "0000000010001000", "1111111110011000", "1111111110100100", "1111111111100110", "0000000000011010", "1111111111111000", "0000000000100001", "1111111111110101", "0000000001000010", "1111111111001110", "1111111110110111", "1111111111110001", "0000000000011101", "0000000000001101", "1111111111111011", "1111111111011110", "0000000000110100", "1111111111100101", "0000000000100011", "1111111111001011", "0000000001011111", "1111111111100100", "1111111111111101", "1111111111011100", "1111111111110111", "1111111111100101", "0000000000100000", "0000000000010010", "1111111111111010", "1111111111100100", "1111111111110010", "0000000000000011", "1111111111010011", "0000000000000000", "0000000001000000", "1111111111101101", "1111111111010101", "1111111111011011", "1111111111100110", "0000000000100011", "0000000000001101", "1111111111111101", "1111111111011000", "0000000000001100", "1111111111011111", "1111111110110001", "0000000000101011", "1111111110111100", "1111111111100100", "0000000000100110", "1111111111111101", "1111111111111010", "0000000000110001", "0000000000100010", "1111111111010110", "1111111110111100", "0000000000001001", "1111111111111011", "0000000000100000", "0000000000001010", "1111111111001111", "1111111111101010", "0000000000001101", "0000000000010001", "1111111111111000", "1111111111100000", "0000000000100010", "0000000000000011", "1111111111110010", "0000000000011001", "1111111111111100", "0000000000010001", "0000000000001111", "1111111111011101", "0000000000010100", "1111111111100111", "1111111111111110", "0000000000101000", "1111111111011100", "0000000000110100", "0000000000110110", "0000000000100101", "1111111111111111", "1111111111001001", "1111111110001010", "0000000000010111", "0000000000000111", "0000000000100110", "1111111110110110", "0000000001011101", "0000000000000010", "1111111111011110", "0000000001000011", "0000000000011110", "1111111111001011", "1111111111110011", "0000000000011001", "1111111111010111", "0000000000000001", "0000000000011011", "0000000000001100", "1111111110111100", "0000000001010010", "1111111111100111", "1111111111101000", "1111111111100110", "1111111111110111", "1111111111101011", "1111111111111001", "0000000000000111", "1111111111100110", "1111111111011111", "1111111111111111", "1111111111110011", "0000000000001001", "0000000000111001", "0000000000001110", "1111111111111110", "0000000000011001", "0000000000101010", "0000000001001110", "1111111110011110", "1111111111101100", "1111111110111100", "0000000010000000", "1111111110100111", "0000000010001011", "1111111111010000", "0000000000001011", "0000000001111001", "0000000000100010", "1111111111011001", "0000000000001111", "1111111101110011", "0000000001100100", "1111111111100111", "0000000001110001", "1111111111001010", "1111111111101010", "0000000001000011", "1111111110110101", "1111111110000100", "0000000001001000", "1111111111010100", "1111111111110101", "1111111111111010", "0000000000011000", "1111111111101001", "0000000000001010", "1111111111010110", "1111111111011001", "0000000000101010", "1111111111011100", "0000000000101000", "1111111111110010", "0000000000000111", "0000000000111000", "0000000000100100", "0000000000011000", "1111111111101001", "0000000000011110", "1111111111010000", "1111111111111111", "1111111111110001", "0000000000001000", "1111111111010100", "1111111111001100", "1111111111001100", "1111111111111110", "1111111111110011", "1111111111011110", "0000000000110010", "1111111111110101", "1111111111100111", "0000000001011101", "0000000000100111", "1111111111110100", "1111111111010011", "1111111111001111", "0000000001011011", "1111111101111100", "0000000000011100", "1111111110110000", "0000000001001010", "0000000000011110", "0000000001000000", "1111111111101111", "0000000000111011", "1111111111100100", "1111111111110101", "0000000000000010", "1111111110100011", "1111111111011100", "0000000001000111", "0000000000100010", "0000000001000111", "1111111111011101", "1111111110111101", "1111111101010010", "1111111111110001", "0000000000101101", "0000000001111101", "0000000000010111", "0000000000011110", "1111111111000010", "0000000000010100", "0000000001000011", "0000000000001110", "1111111110111110", "1111111110010100", "0000000010001010", "0000000000000011", "0000000000000100", "1111111111011110", "1111111111111101", "0000000000001100", "1111111110111100", "0000000001001100", "0000000000100100", "0000000001010110", "1111111111000100", "1111111111110100", "1111111101101100", "0000000000111001", "0000000000010100", "0000000000110011", "1111111111001100", "0000000000110111", "1111111111110110", "0000000000001111", "1111111111010011", "1111111111000100", "1111111111011110", "0000000000110110", "1111111110101110", "1111111111101111", "1111111111101100", "0000000000010111", "0000000000010100", "0000000000111101", "1111111111100011", "1111111110110001", "0000000001100100", "1111111111101001", "1111111110010011", "0000000000000001", "1111111111101111", "1111111111101110", "0000000000010110", "0000000001011101", "1111111110100000", "1111111111111000", "0000000000100101", "1111111111101111", "1111111111000010", "1111111111010010", "0000000000100101", "0000000000101110", "0000000000100111", "0000000001011011", "1111111110111000", "1111111111010101", "0000000001001110", "0000000000000000", "1111111111110110", "0000000000011011", "0000000000001000", "0000000000101010", "1111111111011101", "0000000000011101", "0000000000010000", "1111111111110111", "1111111111101101", "1111111111100101", "1111111111101101", "1111111111101101", "1111111111100001", "0000000000111000", "0000000000001011", "0000000000001111", "0000000001001110", "0000000000000101", "1111111110101000", "0000000001011000", "0000000000000011", "1111111111000000", "0000000000100100", "0000000000000000", "1111111111111011", "1111111111110101", "1111111111001000", "0000000000100101", "0000000000010001", "0000000000011111", "1111111111001110", "1111111111001000", "1111111111000101", "0000000000101010", "1111111111101001", "0000000000011100", "1111111111010010", "0000000001111110", "1111111111111111", "0000000000110010", "0000000001000010", "1111111111100111", "1111111111111010", "0000000000010110", "0000000000010101", "0000000000000111", "0000000000100110", "1111111111100111", "1111111110011110", "0000000000000001", "0000000001010000", "0000000001111001", "1111111111110010", "1111111111000110", "1111111110101111", "1111111111110000", "0000000001011010", "1111111110110011", "1111111110100110", "1111111111101001", "1111111110111100", "1111111111100101", "0000000001000101", "0000000000000000", "0000000000101011", "1111111111100101", "0000000000000000", "0000000000010010", "0000000001010010", "0000000000010010", "1111111111111111", "1111111111011000", "0000000001001011", "1111111111000110", "1111111111000001", "1111111111111010", "1111111110101111", "0000000000100010", "0000000000101101", "0000000001000010", "1111111111110101", "0000000000110101", "0000000000111101", "1111111111000000", "0000000000100011", "1111111111110000", "0000000000000100", "1111111111101010", "0000000000011001", "1111111110111111", "1111111111101011", "1111111111010001", "0000000000101001", "0000000001001001", "0000000000101100", "0000000000000000", "0000000000011100", "1111111111011101", "0000000000101000", "1111111110110000", "1111111111101000", "1111111111001011", "1111111111011001", "0000000000010111", "1111111111111101", "1111111111000111", "1111111111100011", "0000000000011111", "0000000010000001", "0000000000101001", "1111111111001100", "1111111111111011", "0000000000010001", "0000000000011001", "1111111111111001", "1111111111100111", "1111111111111111", "0000000001000110", "0000000000001000", "1111111111110001", "1111111111110011", "1111111111100001", "0000000000000001", "1111111111100000", "1111111111110110", "0000000000000000", "0000000000011110", "0000000000110001", "0000000000011100", "1111111111100110", "1111111111010000", "0000000000000110", "0000000000100100", "0000000001001100", "0000000000111000", "1111111111011001", "1111111111010010", "1111111110111110", "0000000000001111", "1111111111101011", "0000000000010001", "1111111111100111", "1111111111011000", "0000000000101001", "0000000000001110", "1111111111001100", "0000000000000001", "1111111111010001", "1111111111101111", "0000000000000000", "0000000000001011", "0000000000101001", "1111111111111110", "1111111110111001", "0000000000010111", "1111111111101001", "0000000000010101", "0000000000010010", "1111111111011010", "0000000000010100", "0000000000011011", "1111111111111110", "0000000000001100", "1111111111111010", "1111111111100111", "0000000000010111", "1111111111111010", "1111111111011011", "0000000000001101", "0000000000011110", "1111111111001010", "1111111111110100", "0000000000001010", "1111111111101000", "1111111111100110", "0000000001000110", "0000000000000100", "1111111111101001", "1111111111100111", "1111111111111101", "0000000000111101", "1111111111111010", "1111111111011010", "1111111111111010", "0000000000011001", "1111111111001110", "0000000000010101", "0000000000000111", "0000000000010000", "1111111111100111", "0000000000001011", "1111111111011101", "0000000000011111", "1111111111001000", "0000000000011000", "1111111111000111", "1111111111111001", "0000000000110101", "1111111111100110", "1111111111111000", "0000000000011101", "0000000000100010", "0000000000100111", "1111111111001000", "1111111111110100", "0000000000000000", "0000000001100011", "1111111111100001", "0000000000010110", "1111111111100010", "1111111111011011", "0000000000000001", "1111111111101100", "1111111111101010", "0000000000011010", "1111111111011111", "0000000000100110", "1111111110111001", "1111111111110100", "0000000000010101", "0000000001100001", "1111111111000110", "0000000000000011", "0000000000100010", "1111111111000000", "0000000000000110", "1111111111011000", "0000000001100010", "1111111111111110", "0000000000000010", "1111111101111011", "0000000010000000", "1111111111110011", "0000000000111100", "1111111111101101", "1111111111011010", "1111111110111001", "0000000001110110", "0000000000111100", "1111111111111100", "0000000000000001", "1111111111101111", "1111111110101101", "0000000000010010", "1111111111011010", "1111111111101100", "1111111111000000", "0000000001110111", "1111111111011001", "0000000000001010", "1111111111011111", "0000000001010010", "0000000000100000", "0000000001000100", "0000000000000000", "1111111111011001", "1111111111000111", "1111111111101001", "1111111111110001", "0000000000010010", "1111111111110010", "1111111110111111", "0000000000101100", "0000000001000010", "0000000000010010", "1111111111011101", "1111111111101001", "1111111111111000", "0000000001000011", "1111111111100101", "0000000000000000", "1111111110111000", "1111111111010111", "0000000000110001", "0000000000101010", "1111111111101011", "1111111111100100", "1111111111101000", "1111111111111001", "0000000000001110", "0000000000101111", "1111111111000110", "0000000000100111", "0000000000011001", "1111111111101101", "0000000001011000", "1111111110011010", "0000000000000110", "1111111111110011", "0000000000010101", "1111111111100110", "0000000000000011", "0000000000111100", "0000000000001001", "0000000001000110", "0000000000111100", "1111111111110011", "1111111111110110", "1111111111110100", "0000000000010101", "1111111111110110", "0000000000000101", "1111111111001010", "1111111110101011", "0000000000101100", "0000000000110010", "0000000000010001", "1111111110111100", "0000000000010010", "0000000000101001", "0000000000101001", "0000000000010010", "1111111111100111", "1111111111100101", "1111111111111110", "1111111111101011", "0000000000001001", "1111111111110001", "0000000000101110", "0000000000001110", "1111111111010010", "0000000000111100", "0000000000101101", "1111111111101100", "0000000000100111", "1111111111000000", "0000000000100011", "1111111111110100", "1111111111100101", "1111111111000111", "0000000000111011", "1111111111110011", "1111111110110011", "1111111111101101", "0000000000100101", "0000000000100110", "1111111111011100", "0000000001110101", "0000000000001111", "1111111111100100", "0000000000101011", "1111111111110000", "1111111111101010", "1111111111100001", "0000000000001001", "0000000000001100", "1111111111101111", "0000000000010001", "1111111111111011", "0000000000111011", "0000000000100011", "0000000000010011", "1111111111110101", "0000000000000100", "1111111111101100", "0000000000000101", "0000000000101111", "1111111110001010", "0000000000000111", "0000000000000010", "0000000000000111", "0000000000010101", "0000000000010101", "0000000000100010", "1111111111101100", "1111111111110001", "0000000000001000", "1111111111110111", "1111111111100101", "1111111111111000", "1111111111100000", "1111111111001110", "0000000001000001", "0000000000000110", "1111111111011111", "0000000000111101", "1111111111001111", "0000000001110011", "1111111111100110", "1111111111101000", "0000000001001111", "0000000000001001", "1111111111100111", "1111111111100010", "0000000000010011", "0000000000101011", "1111111111011001", "1111111111001111", "0000000000000011", "1111111111001010", "0000000000101010", "0000000000100101", "0000000000000110", "0000000000000011", "1111111111111100", "1111111111111100", "1111111111010100", "1111111111100011", "0000000000111001", "1111111111011000", "1111111111100011", "1111111111100101", "1111111111111110", "1111111111110110", "1111111111110101", "0000000000010101", "1111111111000111", "0000000000010101", "1111111111100000", "0000000000000100", "1111111111100001", "0000000000011111", "0000000000000001", "0000000000100100", "0000000000110111", "0000000001000010", "0000000000110011", "1111111111101000", "1111111111001010", "0000000000000100", "1111111111000110", "1111111111010111", "0000000001110100", "0000000000011001", "0000000000100010", "1111111111111100", "1111111111111011", "0000000000110110", "0000000000100010", "1111111111010000", "1111111111001110", "1111111111111101", "0000000000000000", "1111111111101110", "1111111111000101", "1111111111100000", "0000000000001111", "1111111111100001", "0000000000110000", "0000000000111001", "1111111111010110", "0000000000010011", "0000000000000101", "0000000000000110", "1111111111100000", "1111111111011110", "1111111111110100", "0000000000010000", "1111111111100101", "1111111111101000", "1111111111100000", "0000000000001011", "1111111111010101", "0000000000000000", "0000000000101101", "1111111111111001", "0000000000000111", "1111111111111100", "0000000000000000", "1111111110110111", "1111111111100101", "1111111111000111", "0000000000000111", "0000000000011001", "1111111111010001", "0000000000000011", "0000000001101001", "0000000000001110", "0000000000011011", "1111111110110010", "0000000000111010", "0000000000001101", "1111111111101100", "0000000000101001", "1111111111010100", "0000000000000010", "0000000000011011", "1111111111101110", "1111111111111010", "0000000000001011", "0000000000010101", "0000000000001001", "0000000000101000", "1111111111101010", "1111111111010001", "1111111111010011", "1111111111110011", "1111111111101111", "1111111111110100", "1111111111101111", "0000000000110000", "0000000000001000", "1111111111100011", "1111111111101000", "0000000000000111", "0000000000111011", "1111111111110001", "0000000000100000", "1111111111101100", "1111111111000000", "0000000010110101", "1111111110111111", "0000000010010100", "1111111110011111", "1111111110011010", "0000000011000101", "1111111110111110", "0000000000101011", "0000000000001100", "1111111101000001", "1111111111110110", "0000000001000101", "0000000000100000", "0000000000111001", "1111111101111101", "1111111111011100", "1111111110111001", "0000000000010110", "0000000000000001", "0000000000011011", "1111111110110010", "0000000000101110", "1111111111010100", "0000000000010011", "1111111111110001", "0000000000100010", "1111111111111000", "0000000001000101", "1111111111000001", "0000000000010011", "0000000000101111", "1111111111100111", "1111111111011011", "1111111111101001", "1111111111111011", "0000000000011111", "0000000000001100", "1111111111101001", "1111111111010111", "0000000000010101", "0000000000111001", "1111111111011001", "0000000000001101", "1111111110010101", "0000000000100001", "0000000000100101", "1111111111000001", "1111111110110101", "0000000001101000", "0000000000010110", "1111111111010111", "0000000000001110", "1111111111010011", "0000000000010110", "0000000000000011", "1111111111011001", "0000000000001111", "1111111111000101", "1111111111110110", "0000000000001001", "0000000000101101", "0000000001000011", "1111111111010011", "0000000001100111", "1111111111110110", "1111111111111100", "1111111111100000", "1111111110110010", "1111111110100111", "0000000000000001", "1111111111000101", "0000000000010001", "1111111111111110", "0000000000011110", "1111111111110100", "1111111111011111", "0000000000110100", "1111111111001010", "1111111111001110", "0000000000101001", "1111111110100100", "1111111110100010", "0000000001010011", "1111111111001110", "1111111111100000", "0000000000100010", "1111111111110101", "0000000000100110", "1111111111101001", "0000000001000000", "0000000000100101", "0000000000000011", "1111111111000011", "0000000000010101", "0000000000110111", "0000000000110110", "1111111111100101", "1111111111101110", "0000000000010111", "1111111111110011", "1111111111101010", "0000000000101111", "1111111111110110", "0000000000011100", "0000000001010011", "1111111111100100", "1111111111101110", "1111111110110101", "1111111111100101", "0000000000100000", "1111111111101100", "0000000000011000", "1111111111101010", "0000000000110001", "0000000000001010", "1111111111110011", "0000000000001001", "1111111111111001", "0000000000001100", "1111111111110010", "1111111111000001", "0000000000010110", "1111111111010011", "0000000000110110", "0000000000001010", "0000000000011110", "1111111111011001", "0000000000011111", "0000000000011100", "0000000000000100", "1111111111011110", "1111111111111101", "1111111111011000", "0000000001000011", "0000000000101100", "1111111111110011", "1111111111101011", "1111111111100110", "0000000000110101", "1111111111111111", "1111111111000100", "1111111111111110", "1111111111100100", "0000000001000000", "1111111111111011", "0000000000000011", "1111111111111111", "1111111111100100", "1111111111110101", "1111111111111000", "0000000000001110", "1111111111110000", "0000000000010001", "1111111111110000", "0000000000011111", "1111111111110100", "0000000000110011", "1111111110111100", "0000000000010010", "1111111111111101", "0000000001100001", "1111111110110100", "0000000000110101", "1111111111010101", "0000000000101110", "0000000000011110", "0000000010000010", "1111111111101101", "0000000000101011", "1111111110110001", "0000000000011011", "1111111111000100", "0000000000011011", "0000000000100001", "0000000000110000", "1111111111111000", "0000000000110110", "1111111110101100", "1111111111101110", "1111111111101011", "0000000000001110", "1111111111100111", "0000000000000000", "1111111111110010", "0000000000001111", "1111111111100100", "0000000000000110", "0000000000011010", "1111111111100001", "0000000000001001", "0000000000001001", "0000000000000000", "0000000000010101", "1111111111001011", "1111111111111111", "1111111111101011", "1111111111101011", "1111111111001111", "1111111111101100", "0000000000110011", "0000000000010000", "1111111111010001", "0000000000110001", "1111111110100110", "0000000000011111", "0000000000011101", "0000000000101011", "0000000001101000", "1111111111101011", "1111111111011101", "1111111111001011", "0000000100101111", "1111111111010010", "1111111111100011", "1111111111000010", "1111111111110100", "1111111110000111", "0000000000011011", "1111111111011111", "1111111111101001", "1111111111000100", "0000000000100001", "1111111111111000", "0000000000110100", "0000000000011110", "0000000001011010", "1111111101101101", "1111111111101101", "1111111111100100", "0000000000000101", "1111111111010101", "0000000000101111", "0000000000000101", "1111111111001101", "1111111111110100", "1111111111101100", "0000000000000010", "0000000001011010", "0000000000011010", "0000000000010001", "1111111111101001", "1111111110010100", "0000000000010000", "0000000000011000", "1111111111011100", "1111111110111100", "0000000001011100", "1111111111010110", "0000000000011110", "0000000000101000", "1111111111010101", "0000000000000111", "1111111111010111", "1111111111100000", "1111111111100110", "0000000000100110", "1111111111111101", "1111111111110000", "0000000000001110", "0000000000000101", "0000000000001100", "1111111111111010", "0000000000011111", "0000000000101000", "1111111111010001", "0000000000110101", "1111111111011101", "1111111111000010", "0000000000011110", "0000000000001011", "1111111111011000", "1111111111011011", "1111111111100111", "0000000001000100", "0000000000001101", "0000000000111101", "1111111111000101", "1111111111101011", "0000000000111100", "0000000000101001", "0000000001101000", "1111111111100111", "1111111110100111", "0000000001100011", "1111111110111011", "1111111111100001", "1111111111010101", "0000000000010100", "1111111111110111", "0000000001000111", "0000000000100011", "0000000001001001", "1111111110000101", "0000000000110001", "1111111111101110", "1111111110110101", "0000000000110011", "0000000001001010", "1111111111110010", "1111111110101110", "0000000000011100", "1111111111111110", "1111111111001011", "0000000000101110", "1111111111110101", "1111111111111110", "0000000000000000", "0000000000101111", "1111111111001110", "1111111111110111", "1111111111100110", "1111111111100111", "1111111111010111", "0000000000000010", "0000000000111110", "1111111111100010", "0000000000011110", "1111111111011101", "1111111111100011", "0000000001010100", "0000000000010101", "1111111111000101", "1111111111101110", "0000000000001000", "0000000000000000", "0000000001010001", "0000000001010000", "0000000000010101", "1111111111011101", "1111111111100100", "0000000000000100", "1111111111111100", "0000000001010111", "0000000000010010", "1111111111011001", "0000000001011010", "1111111101101111", "0000000000000000", "0000000000100010", "1111111110001111", "1111111111110100", "0000000000101101", "1111111110011000", "0000000000010001", "1111111111110000", "0000000000001010", "1111111111101001", "0000000001000110", "1111111111111111", "0000000000010101", "1111111111111000", "0000000000000111", "1111111111111011", "0000000000011110", "1111111111011100", "1111111111100001", "1111111110110110", "1111111110111001", "0000000000000000", "0000000000100010", "1111111111100000", "1111111111001100", "0000000001101010", "1111111111111110", "0000000000001001", "1111111111100000", "1111111111111001", "1111111111111110", "0000000000101110", "1111111111010111", "1111111111010110", "0000000000111101", "0000000000010110", "1111111111100111", "0000000000000000", "0000000000001110", "1111111111110011", "0000000000011110", "0000000001000101", "1111111111110011", "0000000000000111", "0000000000001011", "1111111111111000", "0000000001000100", "1111111111110001", "0000000000010001", "1111111110001101", "0000000000010010", "1111111111101100", "0000000001000101", "1111111111010100", "1111111111010011", "0000000000101011", "0000000000110011", "1111111111101011", "1111111111101011", "1111111110100111", "0000000000101110", "0000000001000001", "0000000000100111", "1111111111000101", "1111111110001000", "0000000010000101", "1111111110100111", "1111111111100011", "1111111110110010", "1111111111100011", "0000000000110000", "0000000000110101", "0000000000110010", "1111111111100101", "1111111110111100", "0000000000001101", "1111111111100000", "1111111111100001", "1111111110111100", "0000000001111110", "0000000000011011", "0000000000000100", "1111111111000001", "0000000000110011", "1111111111001110", "0000000000100100", "0000000000011010", "0000000000101000", "0000000000011000", "1111111111101111", "0000000000000000", "1111111111100110", "0000000000000000", "0000000000100001", "0000000000010110", "0000000000001110", "0000000000011111", "1111111111101101", "1111111111100111", "1111111111110001", "1111111111101110", "1111111111110110", "0000000000000110", "1111111111110110", "1111111111011011", "1111111111111000", "0000000000001101", "0000000000101001", "0000000000000001", "1111111111110001", "0000000000000011", "0000000000101110", "1111111111111110", "0000000000000111", "0000000000000001", "1111111111110011", "0000000000011111", "0000000001000001", "1111111111011100", "1111111110101110", "0000000000101011", "1111111111101001", "0000000000011011", "0000000000001111", "0000000000011111", "1111111111110111", "0000000000000111", "0000000000010110", "1111111111010010", "0000000000000001", "0000000000010001", "1111111111111101", "0000000000001100", "1111111111111011", "0000000001010000", "0000000000000100", "0000000000001001", "0000000001000101", "1111111110010011", "0000000001001101", "1111111111000010", "0000000000000100", "1111111111101101", "0000000000101110", "0000000000001101", "0000000000100101", "1111111110110001", "0000000000111010", "1111111111100110", "0000000000100000", "0000000000000000", "0000000000100000", "0000000000011001", "0000000000011100", "1111111110111111", "0000000001010010", "1111111111010011", "0000000000000101", "1111111110011000", "1111111111110111", "1111111111100000", "0000000000000000", "1111111111100110", "1111111111101001", "1111111110110100", "1111111111111100", "1111111110101011", "0000000001101101", "0000000000001111", "0000000000001010", "1111111111100010", "0000000001101001", "1111111111000100", "0000000001100010", "1111111111101101", "1111111111001010", "1111111110101100", "1111111111100011", "1111111111000000", "1111111111100100", "0000000000110011", "0000000000111110", "0000000000111100", "1111111111100000", "0000000000000000", "1111111110110011", "0000000001010100", "1111111111010000", "0000000000110101", "0000000001000100", "1111111110110111", "0000000001011000", "0000000000100000", "1111111110010100", "0000000000000010", "0000000000011001", "0000000000001000", "0000000000000101", "1111111111111101", "0000000000001000", "0000000000110011", "1111111111110000", "1111111111011100", "1111111110101110", "0000000000011011", "0000000000111110", "1111111111001101", "0000000000011100", "0000000000011011", "1111111111111001", "0000000001010110", "0000000000000111", "0000000000010000", "1111111101100001", "0000000000000000", "0000000000011111", "1111111110111101", "1111111111100000", "0000000010111000", "0000000000011010", "1111111111011110", "0000000000111110", "1111111111001001", "1111111111110110", "0000000000100110", "1111111111110000", "0000000010000011", "0000000000010101", "0000000000001010", "1111111110000100", "1111111111110101", "0000000000000001", "1111111111100101", "0000000001111001", "0000000000110001", "0000000000001001", "1111111110110010", "0000000000011111", "1111111101111110", "1111111111010100", "0000000000000110", "1111111110010110", "0000000000101101", "0000000001000001", "1111111111110100", "1111111111011011", "1111111111000111", "1111111110111010", "0000000000000101", "0000000000101011", "0000000000001101", "0000000000100110", "0000000000000000", "1111111111101001", "0000000000011100", "1111111111111001", "0000000000101100", "1111111111001000", "0000000001100110", "1111111111010001", "1111111111101001", "0000000001001110", "1111111111011110", "1111111111000110", "0000000000000110", "1111111111110011", "0000000000100111", "0000000000000111", "0000000000101010", "1111111111010000", "1111111111100000", "0000000000011111", "1111111111111001", "0000000000000000", "0000000000100010", "1111111111000010", "0000000000110011", "0000000000001101", "1111111111011000", "1111111111100111", "0000000001011111", "1111111111000011", "0000000000010100", "0000000000010101", "0000000000010100", "0000000000001011", "1111111111110011", "1111111111010100", "1111111111101010", "0000000000011011", "0000000001000011", "1111111111011000", "1111111111011110", "1111111111100010", "1111111111111000", "1111111110100110", "0000000000101010", "0000000000011101", "1111111111110001", "0000000000101011", "1111111111101010", "1111111111010100", "0000000000011011", "1111111111101110", "1111111111100010", "0000000000010010", "0000000000101101", "1111111110111010", "1111111111001110", "1111111111111101", "0000000001110100", "1111111111111101", "1111111111000111", "1111111111000011", "0000000000101001", "1111111111001000", "0000000001000110", "0000000000000111", "0000000000010000", "1111111111011110", "0000000010100101", "1111111110111000", "0000000001000011", "1111111111101001", "0000000000100010", "1111111111010000", "0000000000011010", "1111111111111001", "0000000000001011", "0000000000111010", "0000000000101001", "1111111111011001", "0000000000010001", "1111111111110110", "0000000000100110", "0000000000010011", "0000000000011011", "1111111111010100", "1111111111111000", "1111111111111100", "0000000000001001", "1111111111011000", "0000000000100111", "0000000001100001", "0000000000101100", "1111111111011111", "1111111101101101", "1111111111011100", "1111111111111101", "0000000000101111", "1111111110001101", "0000000001011111", "1111111111110101", "0000000001011011", "0000000000101110", "1111111111011001", "1111111111010100", "0000000000101100", "0000000001000000", "1111111111001000", "1111111110011111", "1111111111111110", "0000000000001111", "0000000001110000", "0000000001001100", "1111111110111110", "1111111111110110", "1111111111110100", "0000000001010110", "1111111110100011", "1111111110011010", "1111111110110110", "1111111111111101", "1111111110111010", "1111111111000101", "1111111111100011", "1111111111111101", "0000000000001011", "1111111111110000", "0000000000010000", "1111111111110110", "0000000000010001", "1111111111111010", "1111111111011111", "1111111110011011", "0000000000000000", "1111111110001101", "0000000000111101", "0000000000010011", "1111111111101101", "0000000000100111", "0000000000101111", "0000000010001000", "0000000000010111", "1111111111100011", "0000000000000000", "1111111111001001", "0000000000011010", "0000000000100110", "1111111110100000", "1111111111011010", "0000000001000001", "1111111111101000", "1111111111001011", "0000000000011001", "0000000000101000", "0000000000000000", "0000000000001101", "0000000000000111", "1111111111110101", "1111111110111110", "0000000000111100", "1111111111101001", "1111111111110110", "1111111111011110", "0000000000011001", "0000000000011011", "1111111111111101", "0000000000001100", "1111111111011011", "1111111111110100", "1111111111101111", "1111111111111000", "0000000000001010", "1111111111101101", "0000000000000101", "1111111111111001", "0000000000010000", "1111111111111101", "0000000000100010", "0000000000110001", "1111111111011001", "1111111111110011", "0000000000001010", "0000000000010110", "1111111111110100", "0000000000010000", "0000000000001011", "1111111111111001", "0000000000110010", "0000000000100100", "0000000000010111", "1111111111011110", "1111111111110000", "1111111111110110", "0000000000011111", "0000000000001010", "1111111111010010", "1111111111110111", "1111111111110110", "0000000000010110", "1111111111011101", "1111111111010110", "1111111111101111", "0000000000100110", "1111111110110011", "0000000000000000", "0000000000101110", "0000000000001010", "0000000000101010", "1111111111101010", "0000000000101110", "1111111111011001", "1111111110110010", "0000000001110010", "1111111110000111", "0000000001010100", "0000000000110111", "1111111110101110", "0000000000100011", "1111111111111100", "1111111111101000", "0000000000101101", "1111111111010110", "0000000000001001", "1111111111000101", "1111111111011110", "0000000000000000", "1111111111101010", "0000000000001001", "0000000000010110", "1111111111010110", "0000000000111110", "0000000000100001", "1111111111011010", "1111111111110001", "0000000000010000", "0000000000010101", "1111111111111101", "1111111111111001", "0000000000100010", "0000000000001110", "1111111111011010", "1111111111001111", "0000000000011101", "0000000000010110", "0000000000101010", "1111111111100101", "1111111111100011", "1111111111100010", "1111111111010110", "1111111111010010", "0000000000000000", "0000000001000000", "1111111111110010", "0000000000100000", "0000000000100101", "0000000000010000", "0000000000010110", "0000000001100010", "0000000000010100", "1111111110110101", "1111111111111110", "0000000000011111", "1111111111101011", "1111111111110011", "1111111110111101", "0000000001001011", "1111111111110111", "1111111111100001", "0000000001001101", "0000000000011011", "1111111111111101", "1111111111100011", "1111111111001111", "0000000000010000", "0000000000100100", "1111111111110110", "0000000000010001", "1111111111100010", "1111111111111101", "0000000000100001", "1111111111010100", "1111111111110110", "0000000001010110", "0000000000000100", "1111111111101011", "0000000000001110", "1111111111110010", "0000000001001010", "1111111111100101", "1111111111101001", "1111111111100000", "0000000010011111", "1111111111111011", "1111111111101100", "1111111111001101", "1111111111011011", "0000000000010100", "0000000000110001", "0000000000001111", "1111111110111010", "1111111111000100", "1111111111001100", "1111111110101101", "0000000000110001", "0000000000001100", "0000000000010110", "0000000000011111", "1111111111110011", "0000000000100001", "0000000000111000", "1111111111111001", "1111111111110110", "0000000000011011", "0000000000001100", "1111111111111100", "0000000000011110", "1111111111100010", "0000000000011000", "0000000000110011", "0000000000010001", "0000000000000101", "0000000000000100", "1111111110111001", "0000000000001001", "0000000000000001", "0000000001011010", "1111111111110000", "1111111111011000", "1111111111011000", "1111111111101110", "1111111111011100", "1111111111111011", "1111111110110000", "1111111111101101", "1111111111110110", "0000000000111011", "0000000000010110", "1111111111011100", "1111111111100100", "0000000001000001", "0000000000000100", "0000000000010101", "0000000000001010", "1111111111101110", "0000000000011010", "1111111111111101", "1111111111011101", "1111111111100011", "1111111111100101", "0000000000101011", "0000000000010110", "1111111111111001", "0000000000000111", "0000000000000011", "0000000000011101", "1111111111100110", "0000000000010001", "0000000000011101", "1111111111111110", "0000000000000000", "1111111111111100", "0000000000000011", "0000000000000001", "1111111111001111", "1111111111011110", "0000000000010010", "0000000000010011", "0000000000011001", "1111111111010110", "0000000000000010", "1111111111001111", "0000000000000111", "0000000001000000", "0000000001100010", "1111111111101011", "1111111111110101", "0000000001000010", "0000000000001100", "1111111110011001", "0000000000010110", "1111111110110000", "1111111110100100", "0000000001001001", "0000000000110110", "0000000000011101", "1111111111101001", "0000000000010000", "1111111110100101", "0000000001011000", "0000000000001010", "1111111111100110", "1111111111101110", "1111111111101100", "1111111111110010", "1111111111111100", "0000000000011101", "0000000000000111", "1111111111111011", "0000000000101000", "1111111111001111", "0000000000000000", "0000000001000111", "1111111111001101", "0000000000100100", "0000000000000110", "0000000000000011", "1111111110011010", "1111111111111110", "1111111110100101", "0000000000110111", "0000000001000101", "0000000000110100", "1111111110100101", "1111111111110001", "1111111110111101", "0000000000001110", "1111111111110101", "0000000000000001", "1111111110100110", "0000000001011111", "1111111111000010", "1111111111010000", "1111111110011010", "0000000001100100", "0000000000010000", "0000000000011000", "0000000000001000", "1111111111000001", "0000000000101001", "1111111111010110", "0000000001010001", "0000000000011000", "0000000000011110", "0000000000000000", "0000000000000111", "1111111111000011", "0000000000000110", "1111111111101000", "0000000000000111", "1111111111100101", "0000000000011001", "1111111111111101", "1111111111110001", "1111111111101110", "0000000000110111", "1111111111011111", "1111111111010000", "0000000001011011", "0000000000011110", "0000000000011111", "1111111111110101", "0000000000011101", "1111111111001011", "1111111111111011", "1111111111111100", "1111111111111111", "1111111110110000", "1111111111111001", "0000000000011010", "0000000001100110", "1111111111010101", "0000000000000000", "1111111110111001", "1111111111011101", "1111111111110010", "0000000000101100", "1111111111110000", "1111111111011101", "0000000001010100", "1111111111101111", "0000000000010101", "1111111111101001", "1111111111110101", "1111111111100110", "0000000000010000", "0000000000001000", "1111111111110000", "0000000000101100", "0000000000011100", "0000000000011011", "0000000000000100", "1111111111110000", "1111111111101000", "0000000000001011", "1111111111111101", "0000000000010100", "1111111111100100", "0000000000000000", "0000000000001001", "0000000000001101", "0000000000011001", "1111111111010100", "1111111111100111", "1111111111010110", "0000000000011101", "1111111111110100", "1111111111010110", "1111111111101110", "0000000000100101", "0000000000010011", "1111111111101101", "1111111111111111", "1111111111011101", "0000000000010101", "0000000000011101", "0000000000100001", "1111111111100011", "0000000000101010", "1111111111111000", "1111111111110010", "0000000000010101", "0000000000000001", "1111111111100100", "0000000000011011", "0000000000100100", "1111111111101011", "0000000000100010", "0000000000100110", "1111111111011110", "1111111111011110", "0000000000011001", "1111111110111010", "1111111111000101", "1111111111111011", "1111111111111010", "1111111111011100", "0000000000001111", "1111111110111011", "0000000011000101", "0000000000101011", "0000000000000000", "1111111110110011", "0000000000001101", "1111111111100001", "0000000000010001", "1111111111100001", "1111111111001111", "1111111111111111", "1111111111001101", "0000000010001001", "0000000000101011", "0000000000110110", "1111111111101100", "1111111101111000", "0000000000110110", "0000000000111101", "1111111111000101", "0000000001000100", "1111111111010001", "1111111111001001", "0000000000010011", "0000000000001000", "0000000000001101", "1111111110111110", "0000000000010110", "0000000000001110", "0000000000011001", "0000000000000100", "0000000000000011", "0000000000111000", "0000000000010111", "1111111111010001", "1111111111101001", "1111111111111111", "0000000000011001", "0000000000110101", "1111111111100000", "0000000000000011", "0000000000000000", "0000000000011101", "0000000000100011", "1111111111110100", "1111111111011100", "0000000000011000", "1111111111011100", "0000000000110001", "0000000000001100", "0000000001000111", "0000000000000010", "1111111111010010", "0000000001000110", "0000000010011101", "1111111111111000", "1111111111101110", "1111111101000101", "0000000001111111", "0000000010000110", "0000000000111000", "1111111111010100", "1111111110010100", "1111111101010100", "1111111110100000", "0000000001000110", "0000000001010011", "1111111110111000", "0000000000011100", "0000000001000100", "0000000000110110", "0000000000101100", "0000000000000111", "1111111110101111", "0000000000000000", "1111111111000111", "0000000000000101", "0000000001100111", "0000000001111111", "1111111110101010", "1111111111000000", "1111111111111101", "1111111111110010", "0000000000000101", "0000000000000111", "1111111111000100", "0000000001010101", "1111111111100010", "0000000000000110", "1111111110101001", "0000000000101110", "0000000000111001", "1111111111000010", "0000000000110001", "1111111110111010", "0000000000011000", "0000000001010111", "1111111110000001", "1111111111111111", "1111111110111011", "0000000001001011", "0000000001111110", "0000000000101110", "1111111110111000", "1111111111110000", "0000000000010000", "0000000001101000", "1111111111010110", "0000000000010000", "1111111111010110", "0000000000010001", "0000000001001000", "0000000000010001", "1111111111100110", "0000000000001000", "1111111111111100", "1111111111101010", "1111111111110110", "0000000000001001", "1111111111110001", "1111111111100100", "1111111110111111", "0000000000011010", "0000000000101100", "0000000001000000", "0000000001001010", "0000000000111000", "1111111111011011", "1111111111011111", "1111111110101011", "0000000000011101", "1111111111111110", "1111111111111100", "0000000000100000", "1111111111111101", "0000000000100100", "0000000000111111", "1111111111001101", "1111111111010010", "0000000000000110", "0000000000010001", "0000000000100110", "1111111111001110", "0000000000001001", "1111111111100010", "1111111111111000", "0000000000000001", "0000000000001100", "1111111111010011", "1111111111111010", "1111111111110110", "0000000000000010", "1111111111011111", "0000000000001001", "1111111111011100", "1111111111101000", "0000000000001010", "1111111111110000", "1111111110010011", "0000000001011000", "1111111110110110", "0000000010100111", "0000000000111111", "1111111111101100", "1111111110110110", "0000000000010110", "1111111110110001", "0000000000001000", "0000000000000000", "1111111111101101", "1111111111110110", "0000000000011001", "1111111111110110", "0000000001000100", "0000000000011001", "1111111111110000", "1111111110000011", "1111111111110011", "0000000000000110", "1111111111110101", "0000000000010011", "0000000000001100", "0000000000101100", "0000000000000010", "0000000000000100", "1111111111000110", "0000000000101000", "1111111111000011", "0000000000011001", "0000000000110110", "0000000001001001", "1111111111011101", "0000000001011001", "1111111111001101", "1111111100111110", "0000000000001101", "0000000001000011", "0000000000110110", "1111111111100111", "0000000000100000", "0000000000101010", "0000000010100101", "1111111111101010", "1111111111110111", "1111111111111110", "0000000000101110", "1111111111000101", "0000000000101111", "1111111110110110", "0000000010010011", "1111111111101000", "1111111110111111", "1111111110110111", "1111111111011100", "0000000001010101", "0000000000000110", "1111111111100010", "1111111111101001", "0000000001000110", "0000000000101111", "1111111111110001", "1111111111011000", "0000000000000000", "1111111111011100", "1111111111010011", "1111111111100010", "0000000001001100", "1111111111110011", "0000000000101010", "0000000000011010", "0000000000110101", "0000000000101011", "1111111111001011", "1111111111010010", "0000000000011100", "1111111111111101", "0000000000001000", "0000000000101001", "0000000010000001", "1111111111101101", "1111111111100010", "1111111110000101", "1111111111100001", "0000000000010110", "1111111111110001", "1111111111011101", "0000000001011011", "1111111111100111", "0000000001010001", "1111111110110101", "1111111110111010", "0000000000010001", "1111111110111000", "0000000000001110", "1111111111110110", "1111111111110101", "0000000010111111", "1111111110000100", "1111111111010011", "1111111110011000", "0000000000101101", "0000000001001011", "0000000001000000", "1111111111111000", "0000000000000000", "1111111111101110", "0000000000101011", "1111111110111111", "1111111110100000", "1111111111100000", "0000000000110011", "0000000000111110", "1111111111101110", "1111111111111010", "0000000000010011", "0000000000000001", "1111111111110000", "0000000000100010", "0000000000010101", "0000000000010100", "1111111111110111", "0000000000001100", "0000000000010110", "1111111111110111", "1111111111111111", "0000000000011110", "0000000000100010", "1111111111101111", "0000000000010110", "1111111111011011", "0000000001000101", "0000000000010111", "1111111111100110", "1111111111001010", "0000000000000001", "1111111111000110", "0000000001011100", "1111111111010010", "0000000000011100", "1111111111001100", "0000000000000001", "1111111111101100", "0000000000001110", "1111111111011101", "0000000000011010", "1111111111011011", "0000000000010000", "0000000000000101", "1111111110111001", "1111111111111001", "0000000000100010", "0000000000111001", "0000000000000001", "1111111111100001", "1111111111001101", "0000000001000100", "1111111110110110", "0000000001000100", "0000000000010100", "1111111111001001", "0000000001001100", "1111111111111010", "0000000000001010", "1111111110000101", "1111111110111100", "0000000000010110", "1111111111001101", "0000000000101001", "0000000010000100", "1111111111101110", "0000000010010101", "1111111111011000", "1111111111111000", "1111111110101011", "0000000000000011", "1111111111000010", "0000000000011011", "1111111111101110", "0000000000000011", "0000000000010000", "0000000000000010", "1111111111001110", "0000000000011011", "0000000000101110", "0000000000001111", "0000000000010110", "1111111111110000", "1111111111101110", "0000000000000100", "1111111111100110", "0000000000000000", "0000000000000000", "1111111111100100", "1111111111110110", "1111111111100011", "0000000000101110", "1111111111100110", "0000000010001110", "0000000010010001", "1111111101111011", "0000000000111110", "1111111110100001", "1111111110011001", "1111111111100111", "1111111111000100", "0000000000001100", "1111111110010000", "0000000000010011", "0000000001110001", "1111111111010111", "0000000000001010", "0000000000110001", "0000000000001010", "1111111111110111", "1111111111010100", "1111111111011101", "0000000000101010", "1111111111010100", "0000000001011001", "1111111111010101", "0000000000011011", "1111111111011000", "1111111111110100", "1111111111111111", "0000000000000101", "0000000000001101", "1111111111110101", "0000000000100001", "1111111111111010", "1111111111111000", "0000000000101101", "1111111111111110", "0000000000000110", "1111111111100000", "0000000000100100", "1111111111111000", "0000000000001011", "1111111111110001", "1111111101010101", "0000000000010011", "0000000000000101", "0000000001101000", "1111111111000101", "0000000001100001", "0000000000001100", "1111111111100000", "1111111111111011", "1111111110100001", "1111111110001001", "1111111110111010", "0000000000011111", "0000000001101001", "0000000000101101", "0000000001010100", "1111111110000010", "1111111111100111", "0000000000110011", "1111111111011000", "0000000000000111", "0000000001110110", "1111111111101011", "1111111111010100", "0000000000011010", "1111111111010101", "1111111111010100", "0000000000010101", "1111111111101011", "0000000000011011", "1111111111111010", "1111111111101111", "0000000000011000", "0000000000011011", "0000000000011110", "1111111111011001", "0000000000000000", "0000000000001111", "1111111111101100", "1111111111100110", "0000000000000100", "1111111111101101", "0000000000101011", "0000000001001001", "0000000000000110", "0000000000000100", "1111111110110011", "0000000000001000", "1111111111111101", "0000000000000000", "1111111110001101", "0000000000111011", "1111111111111110", "0000000000010111", "0000000000011000", "1111111111001111", "1111111110100010", "1111111111010110", "0000000000001111", "0000000001101100", "1111111111000110", "0000000000110101", "1111111111100010", "0000000000100101", "0000000000100011", "1111111111110100", "0000000000001000", "1111111111011011", "1111111111101000", "1111111111110111", "1111111111100100", "1111111111100111", "0000000000011111", "0000000000010101", "0000000000011111", "0000000000010111");
    Plus214_i_1 <= ("1111111111110011", "0000000000010101", "1111111111110100", "1111111111110010", "0000000000100011", "1111111111100000", "0000000000000111", "0000000000010001", "0000000000000001", "1111111111110101");
    process(all)
    begin
        next_feedback <= feedback;
        next_state <= state;
        next_was_valid <= was_valid;
        valid_out <= '0';
        output <= (others => (others => '0'));
        Block386_i_0 <= (others => (others => '0'));
        Block386_valid_in <= '0';
        Convolution28_i_0 <= (others => (others => '0'));
        Convolution28_valid_in <= '0';
        Plus30_i_0 <= (others => (others => '0'));
        Plus30_valid_in <= '0';
        ReLU32_i_0 <= (others => (others => '0'));
        ReLU32_valid_in <= '0';
        Pooling66_i_0 <= (others => (others => '0'));
        Pooling66_valid_in <= '0';
        Convolution110_i_0 <= (others => (others => '0'));
        Convolution110_valid_in <= '0';
        Plus112_i_0 <= (others => (others => '0'));
        Plus112_valid_in <= '0';
        ReLU114_i_0 <= (others => (others => '0'));
        ReLU114_valid_in <= '0';
        Pooling160_i_0 <= (others => (others => '0'));
        Pooling160_valid_in <= '0';
        Times212_i_0 <= (others => (others => '0'));
        Times212_valid_in <= '0';
        Plus214_i_0 <= (others => (others => '0'));
        Plus214_valid_in <= '0';

        case state is
            when 0 =>
                next_state <= 0;
                if valid_in then
                    next_state <= 2;
					next_was_valid <= '1';
                end if;
            when 1 =>
                Block386_i_0 <= input(783 downto 0);
                Block386_valid_in <= '1';
                if Block386_valid_out then
                    next_state <= 2;
                    next_feedback(783 downto 0) <= Block386_o;
                end if;
            when 2 =>
                Convolution28_i_0 <= input(783 downto 0);
                Convolution28_valid_in <= '1';
                if Convolution28_valid_out then
                    next_state <= 3;
                    next_feedback(6271 downto 0) <= Convolution28_o;
                end if;
            when 3 =>
                Plus30_i_0 <= feedback(6271 downto 0);
                Plus30_valid_in <= '1';
                if Plus30_valid_out then
                    next_state <= 4;
                    next_feedback(6271 downto 0) <= Plus30_o;
                end if;
            when 4 =>
                ReLU32_i_0 <= feedback(6271 downto 0);
                ReLU32_valid_in <= '1';
                if ReLU32_valid_out then
                    next_state <= 5;
                    next_feedback(6271 downto 0) <= ReLU32_o;
                end if;
            when 5 =>
                Pooling66_i_0 <= feedback(6271 downto 0);
                Pooling66_valid_in <= '1';
                if Pooling66_valid_out then
                    next_state <= 6;
                    next_feedback(1567 downto 0) <= Pooling66_o;
                end if;
            when 6 =>
                Convolution110_i_0 <= feedback(1567 downto 0);
                Convolution110_valid_in <= '1';
                if Convolution110_valid_out then
                    next_state <= 7;
                    next_feedback(3135 downto 0) <= Convolution110_o;
                end if;
            when 7 =>
                Plus112_i_0 <= feedback(3135 downto 0);
                Plus112_valid_in <= '1';
                if Plus112_valid_out then
                    next_state <= 8;
                    next_feedback(3135 downto 0) <= Plus112_o;
                end if;
            when 8 =>
                ReLU114_i_0 <= feedback(3135 downto 0);
                ReLU114_valid_in <= '1';
                if ReLU114_valid_out then
                    next_state <= 9;
                    next_feedback(3135 downto 0) <= ReLU114_o;
                end if;
            when 9 =>
                Pooling160_i_0 <= feedback(3135 downto 0);
                Pooling160_valid_in <= '1';
                if Pooling160_valid_out then
                    next_state <= 10;
                    next_feedback(255 downto 0) <= Pooling160_o;
                end if;
            when 10 =>
                Times212_i_0 <= feedback(255 downto 0);
                Times212_valid_in <= '1';
                if Times212_valid_out then
                    next_state <= 11;
                    next_feedback(9 downto 0) <= Times212_o;
                end if;
            when others =>
                Plus214_i_0 <= feedback(9 downto 0);
                output(9 downto 0) <= Plus214_o;
                Plus214_valid_in <= '1';
                valid_out <= Plus214_valid_out;
                if not valid_in then
                    next_was_valid <= '0';
                    valid_out <= '0';
                elsif not was_valid then
                    next_was_valid <= '1';
                    next_state <= 0;
                end if;
        end case;
    end process;

    process(clk, rst)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                feedback <= (others => (others => '0'));
                state <= 0;
                was_valid <= '0';
            else
                feedback <= next_feedback;
                state <= next_state;
                was_valid <= next_was_valid;
            end if;
        end if;
    end process;
end Behavioral;
