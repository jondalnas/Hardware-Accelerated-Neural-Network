library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;


use work.types.all;
use work.defs.all;

entity nn_tb is
end nn_tb;

architecture nn_test of nn_tb is
    signal input : array_type(28 * 28 - 1 downto 0)(DATA_WIDTH - 1 downto 0);
    signal output : array_type(10 - 1 downto 0)(DATA_WIDTH - 1 downto 0);
    
	signal clk, rst, valid_in, valid_out : std_logic := '0';
begin
	clk <= not clk after 5 ns;

    nn : entity work.nn
        generic map(
            data_width => DATA_WIDTH,
			num_in => NN_INPUT,
			num_out => NN_OUTPUT,
			num_feedback => NN_FEEDBACK
        )
        port map (
			clk => clk,
			rst => rst,
			valid_in => valid_in,
			valid_out => valid_out,
			input => input,
			output => output
        );
        
        
    process
		constant BLACK : signed := "0000000100000000";
		constant WHITE : signed := "0000000000000000";
		constant GRAYE : signed :=  "0000000010000000";
        variable seed1, seed2 : integer := 999;
        
        impure function rand_slv(len : integer) return std_logic_vector is
            variable r : real;
            variable slv : std_logic_vector(len - 1 downto 0);
        begin
            for i in slv'range loop
                uniform(seed1, seed2, r);
                if r > 0.5 then 
                    slv(i) := '1';
                else
                    slv(i) := '0';
                end if;
            end loop;
            return slv;
        end function;
    begin
		rst <= '1';
		wait for 200 ns;
		rst <= '0';

            -- 1
            input <= (  X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"000a", X"0015", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"004e", X"00e6", X"00fb", X"0039", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0072", X"0100", X"0100", X"0100", X"006e", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0039", X"0100", X"0100", X"0100", X"0100", X"006e", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0039", X"00cc", X"0100", X"00f0", X"0100", X"0100", X"006e", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"003f", X"0092", X"0100", X"0100", X"0100", X"0073", X"0100", X"0100", X"006e", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"007b", X"0100", X"0100", X"0100", X"00f2", X"0078", X"002e", X"0100", X"0100", X"006e", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0068", X"00fb", X"0100", X"0100", X"009d", X"001f", X"0000", X"0049", X"0100", X"0100", X"0039", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0032", X"00fb", X"0100", X"0100", X"0059", X"0000", X"0000", X"0000", X"0068", X"0100", X"0100", X"001f", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"000a", X"00e5", X"0100", X"00fb", X"0049", X"0000", X"0000", X"0000", X"0000", X"006e", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0010", X"00f2", X"0100", X"007d", X"0000", X"0000", X"0000", X"0000", X"0000", X"006e", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0025", X"003f", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"006e", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0088", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0092", X"0100", X"00db", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0092", X"0100", X"00db", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0092", X"0100", X"00db", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0088", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"006e", X"0100", X"0100", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"006e", X"0100", X"0100", X"0010", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0054", X"0100", X"0100", X"0025", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0049", X"0100", X"0100", X"0025", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"002a", X"0049", X"0020", X"000a", X"0025", X"0010", X"0000", X"002a", X"0049", X"0049", X"0088", X"0100", X"0100", X"0025", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"002a", X"00fb", X"0100", X"0100", X"0100", X"0100", X"0100", X"00e6", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"00e1", X"00db", X"00f6", X"0100", X"0100", X"00e6", X"0063", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"001f", X"00f0", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"0100", X"00d1", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0010", X"0039", X"0069", X"006e", X"0063", X"0083", X"0092", X"007d", X"0034", X"0029", X"0049", X"0068", X"0092", X"0092", X"0092", X"0092", X"006e", X"0078", X"0092", X"002f", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000",
                        X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000", X"0000");

--		input <= (WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, BLACK, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, BLACK, BLACK, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, BLACK, BLACK, BLACK, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, BLACK, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, BLACK, BLACK, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, BLACK, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, GRAYE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE,
--				  WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE, WHITE);

		valid_in <= '1';
        
        wait until valid_out = '1';
        wait for 10 ns;
		valid_in <= '0';

		wait until valid_out = '0';
		wait for 1 ms;
		valid_in <= '1';
		wait for 1 ms;
    end process;
end nn_test;
