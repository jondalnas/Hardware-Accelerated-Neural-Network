library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.types.all;

package defs is
-- INSTRUCTIONS
-- INPUT SIZE
    constant INST_SIZE : Integer := 3;
end defs;
