library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.types.all;
use IEEE.NUMERIC_STD.ALL;

entity nn is
    generic(
        num_in : positive;
        num_out : positive;
        num_feedback : positive;
        data_width : integer
    );
    Port (
        clk : in std_logic;
        rst : in std_logic;
        valid_in : in std_logic;
        valid_out : out std_logic;
        input : in array_type(num_in-1 downto 0);
        output : out array_type(num_out-1 downto 0)
     );
end nn;

architecture Behavioral of nn is
    signal feedback, next_feedback : array_type(num_feedback-1 downto 0);
    signal was_valid, next_was_valid : std_logic;

    constant num_states : positive := 11;
    signal state, next_state : integer;

    signal Block386_o : array_type(783 downto 0)(data_width-1 downto 0);
    signal Block386_i_0 : array_type(783 downto 0)(data_width-1 downto 0);
    signal Block386_i_1 : array_type(0 downto 0)(data_width-1 downto 0);
    signal Convolution28_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Convolution28_i_0 : array_type(783 downto 0)(data_width-1 downto 0);
    signal Convolution28_i_1 : array_type(199 downto 0)(data_width-1 downto 0);
    signal Plus30_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Plus30_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Plus30_i_1 : array_type(7 downto 0)(data_width-1 downto 0);
    signal ReLU32_o : array_type(6271 downto 0)(data_width-1 downto 0);
    signal ReLU32_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Pooling66_o : array_type(1567 downto 0)(data_width-1 downto 0);
    signal Pooling66_i_0 : array_type(6271 downto 0)(data_width-1 downto 0);
    signal Convolution110_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Convolution110_i_0 : array_type(1567 downto 0)(data_width-1 downto 0);
    signal Convolution110_i_1 : array_type(3199 downto 0)(data_width-1 downto 0);
    signal Plus112_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Plus112_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Plus112_i_1 : array_type(15 downto 0)(data_width-1 downto 0);
    signal ReLU114_o : array_type(3135 downto 0)(data_width-1 downto 0);
    signal ReLU114_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Pooling160_o : array_type(255 downto 0)(data_width-1 downto 0);
    signal Pooling160_i_0 : array_type(3135 downto 0)(data_width-1 downto 0);
    signal Times212_o : array_type(9 downto 0)(data_width-1 downto 0);
    signal Times212_i_0 : array_type(255 downto 0)(data_width-1 downto 0);
    signal Times212_i_1 : array_type(2559 downto 0)(data_width-1 downto 0);
    signal Plus214_o : array_type(9 downto 0)(data_width-1 downto 0);
    signal Plus214_i_0 : array_type(9 downto 0)(data_width-1 downto 0);
    signal Plus214_i_1 : array_type(9 downto 0)(data_width-1 downto 0);
begin
    Block386 : entity work.div
        generic map (
            input_size => 784,
            data_width => 16
        )
        port map (
            a => Block386_i_0,
            b => Block386_i_1,
            c => Block386_o
        );
    Convolution28 : entity work.conv
        generic map (
            num_dimensions => 2,
            dimensions_x => (1, 1, 28, 28),
            x_size => 784,
            dimensions_w => (8, 1, 5, 5),
            w_size => 200,
            kernel_shape => (5, 5),
            dilation => (1, 1),
            stride => (1, 1),
            data_width => 16,
            y_size => 6272
        )
        port map (
            x => Convolution28_i_0,
            w => Convolution28_i_1,
            y => Convolution28_o
        );
    Plus30 : entity work.add
        generic map (
            input_size => 6272,
            data_width => 16
        )
        port map (
            a => Plus30_i_0,
            b => Plus30_i_1,
            c => Plus30_o
        );
    ReLU32 : entity work.relu
        generic map (
            input_size => 6272,
            data_width => 16
        )
        port map (
            x => ReLU32_i_0,
            y => ReLU32_o
        );
    Pooling66 : entity work.max_pool
        generic map (
            num_dimensions => 2,
            kernel_shape => (2, 2),
            pads => (0, 0, 0, 0),
            strides => (2, 2),
            in_dimensions => (1, 8, 28, 28),
            input_size => 6272,
            output_size => 1568,
            data_width => 16
        )
        port map (
            x => Pooling66_i_0,
            y => Pooling66_o
        );
    Convolution110 : entity work.conv
        generic map (
            num_dimensions => 2,
            dimensions_x => (1, 8, 14, 14),
            x_size => 1568,
            dimensions_w => (16, 8, 5, 5),
            w_size => 3200,
            kernel_shape => (5, 5),
            dilation => (1, 1),
            stride => (1, 1),
            data_width => 16,
            y_size => 3136
        )
        port map (
            x => Convolution110_i_0,
            w => Convolution110_i_1,
            y => Convolution110_o
        );
    Plus112 : entity work.add
        generic map (
            input_size => 3136,
            data_width => 16
        )
        port map (
            a => Plus112_i_0,
            b => Plus112_i_1,
            c => Plus112_o
        );
    ReLU114 : entity work.relu
        generic map (
            input_size => 3136,
            data_width => 16
        )
        port map (
            x => ReLU114_i_0,
            y => ReLU114_o
        );
    Pooling160 : entity work.max_pool
        generic map (
            num_dimensions => 2,
            kernel_shape => (3, 3),
            pads => (0, 0, 0, 0),
            strides => (3, 3),
            in_dimensions => (1, 16, 14, 14),
            input_size => 3136,
            output_size => 256,
            data_width => 16
        )
        port map (
            x => Pooling160_i_0,
            y => Pooling160_o
        );
    Times212 : entity work.mat_mul
        generic map (
            num_dimensions => 0,
            a_dim => (1, 256),
            b_dim => (256, 10),
            a_size => 256,
            b_size => 2560,
            y_size => 10,
            data_width => 16
        )
        port map (
            a => Times212_i_0,
            b => Times212_i_1,
            y => Times212_o
        );
    Plus214 : entity work.add
        generic map (
            input_size => 10,
            data_width => 16
        )
        port map (
            a => Plus214_i_0,
            b => Plus214_i_1,
            c => Plus214_o
        );

    Block386_i_1 <= (0 => "0111111111111111");
    Convolution28_i_1 <= ("1111111011011101", "1110000110101110", "1011111011011111", "1111011110111101", "0001001000100110", "1011010000111011", "1100001100101010", "1111100110101111", "0110001001010100", "0010000110111001", "1100000100001110", "0000011100011110", "0111111111111111", "0100011100000000", "1100011101111000", "1110101110010101", "0100011101011101", "0100101111001001", "1101101001000110", "1011000110000100", "0000010011101101", "0001110011101110", "1110010000000111", "1100001011101100", "1101101010101010", "1111101011100110", "0001101111111011", "0011111111010110", "0011011000111010", "0000011000110110", "1111001100001101", "1101110010001111", "1111111101110000", "0100001101111010", "0011001110100010", "1110110010110010", "1101011000101111", "1110101110100111", "0010110111110011", "0010111110110010", "1011011101010111", "1100111010100001", "1110100111000101", "0001110100110000", "0010101010010111", "1100111101000011", "1110001010100001", "1111011110000110", "1111111000100011", "0010010001110111", "1111110011111000", "0000110101100000", "0010000001110110", "0010111001001110", "0101100001110001", "0010101011011110", "0011010101100000", "0011000101000010", "0010101000101010", "0001111100011011", "1100001111110110", "1111011001000111", "1110110110000001", "1110100111001001", "1110000001101010", "1000001110000000", "1010010001100111", "1011101100011100", "1011000100001110", "1100011010011010", "1110011010001000", "1101010101010101", "1101001101010010", "1110110101001111", "1111011111011101", "1101101000110010", "1101010101110100", "1101011000000101", "1111010111011101", "1110001110001000", "1100001011111010", "1110010100001000", "1111100010100011", "0001010011110101", "0001010010111011", "1100110111011100", "1111110011111110", "0000111111000111", "0000010101101101", "0001110100110000", "0000110000011001", "0010111110011110", "0001110000010100", "1111111010010001", "0001011100110000", "0010100111101100", "0010110011110001", "0000001110111000", "0001101011000111", "0010101110011100", "1110010010001010", "1111000001100001", "1111111110110010", "1110001100011011", "1110101101011111", "0000101101100101", "0001101000111100", "1110101111111101", "1110001100011110", "1011100000001110", "1111100001001011", "0011010010001001", "1111111000100110", "1100001100110110", "1011011111001110", "1111000100110110", "0001001000110000", "0010001101101100", "0000010101110011", "1111111010000110", "0000000100111101", "0001111110000000", "0101000000010100", "0101011101110101", "0001111000110111", "1110101011000000", "1101010101000110", "1110011110000111", "0000011011011001", "0001001000011111", "0001011101101000", "1011100111011001", "1010001000100100", "1011010010110100", "1100111011010010", "0100010100101000", "0010110001001101", "1101111110110101", "1101001110100101", "1110010100000001", "0001110000101101", "0101010001010111", "0010111010110001", "0001000010001111", "1111000111111010", "0000011110110101", "0010011011000011", "0001111001010101", "0011110000001101", "0001110010010100", "0000110010001010", "0100011110011101", "1110010010001110", "1100010101101011", "1110010011100011", "0010111010100100", "0011111001011000", "1100101111010010", "1100100100010000", "1110000001010001", "0011010100011100", "0010011001100110", "1100010101100100", "1101100100011010", "1111010010001010", "0010001110010111", "0000111010100101", "1110100111110010", "1101001011111101", "1110110010001011", "0010110010100001", "0001011111001000", "0000100100010010", "0001000100101100", "1111101000010111", "1111110100101101", "1110111100011011", "0000101110111100", "0001110110100101", "0010101101111100", "0001010100100000", "0011000000110000", "0001100011110110", "0010100001010111", "0100100010011000", "1111000011100110", "0001100100010101", "0001000011110111", "0000011000011101", "0001000100011011", "0000001110100001", "1110111000110001", "1111000010001011", "1110011010111000", "1011111110110110", "1111101101101011", "1110011110110100", "1100100101000111", "1101101110001110", "1110011110100011");
    Plus30_i_1 <= ("1110101101010011", "1100100001111001", "0000101110111010", "1111110111011000", "1111011110101110", "1110111100100100", "0000001010011101", "1111000010000000");
    Convolution110_i_1 <= ("1111100111001001", "1111010001011010", "1111111100101001", "1110111110010001", "0000110111110000", "0000101011001000", "1110101001110011", "1101110101000110", "1111110110010001", "0000100011011101", "0000010100010110", "1111111001111111", "1111011111101010", "1110110010110001", "1111000110011100", "0000100011110001", "0000000000011001", "0000101010101011", "1110100011010100", "1111000011010101", "0000000001101110", "0010000000101010", "0001100011001000", "1111100100000110", "1110111110011010", "1100100110111001", "1101110101011101", "1101111011001011", "0000101001011111", "0000101101000010", "0000000100111110", "1110001010100011", "1111011111001111", "0000001011001010", "1111100110100110", "0001010110110001", "0001111000101000", "1111110110000100", "1110111010111000", "1111101010000110", "1111011110001100", "0001011111010011", "0001011100111010", "1110110101110101", "0000001111011010", "1110111000011010", "0000111010001010", "0000110101110010", "0000011010010000", "0000011101100101", "1110110000100111", "1110111011011010", "0000101000011000", "0000111011101001", "1110111010101111", "1111000000010000", "1110010101111101", "1110110111000110", "1111100000100011", "1111010100100101", "1110011111000001", "1110001111000011", "1110010001001000", "1111010011101000", "0000100001001110", "1101111011010000", "1111001010110011", "1101010101100010", "1110111011000100", "1111101111110100", "0000001110011110", "0000101101110110", "1111001000010110", "1110100000000010", "1110001101011011", "0000110100110101", "1111100111101001", "1111110010011100", "1111110101000000", "0000001110101100", "0000011000100000", "1111111111001110", "0000110101001011", "1111010010111100", "1111100011111001", "0000100111010001", "0000001101100001", "1101111100000010", "1101101110010110", "1110010101001100", "0000001001001010", "0000100010101101", "1111101110011011", "1101100100000011", "1110111111001011", "1111111010101011", "0000111100000111", "0001010110111110", "1111011101101011", "0000011100001011", "0001011001100001", "1111011110011110", "1110111000110110", "1101100010000000", "1111001010100000", "0000101111010111", "0010011001100101", "0000011111010011", "1110001101011000", "1110010000100010", "1111010011100111", "0000010001101011", "0000111110011000", "1110110110100101", "1110110111101001", "1100100111010011", "1111101101111000", "0000011011001110", "0000001100011000", "1111110111110010", "1111000010010111", "1110101100110000", "1111001110011110", "0000010010010000", "0000000110111011", "0001001001101001", "0000001010000101", "1101010011011000", "1110001101110000", "1110101101000011", "0001010101101111", "0011100111011100", "0010001001000111", "1111000000000110", "1110010000010001", "1110110011101001", "1111011001000101", "0010000011110101", "0000110100101011", "0000100001010100", "1100101000100000", "1101100000100011", "1111101101100100", "0000010111111101", "0000111010101000", "1111100100110000", "1110111010010011", "1101110111101001", "1110010010111011", "1111110000001010", "0000011011110100", "1110101000101101", "1101101011101010", "1111101010110011", "1110000001101111", "0000110010110101", "0001100011111101", "1111001101110000", "1101110101100001", "1110110011010101", "1111010100001100", "0000000001000000", "0000011011101100", "0000010111111011", "1110101101100010", "0000001011111010", "0000100001011001", "0001111101111010", "0000011111000011", "0000000110100100", "1111001111100001", "1111001001110101", "0001110101011011", "0001101000100110", "1111010001111111", "1110000001010001", "0001001001110111", "0000011010100110", "1111110011101111", "0000110011001100", "1111100010110001", "1111011001001011", "1111100010100110", "0000011010001100", "0000101100010101", "0000011111111000", "1110110000111010", "1110111000000100", "0000001010010110", "0000001110001001", "1111001011111110", "0000001110101101", "1110111110011110", "1110001011110010", "1101110110011001", "0001000100001110", "0000100111111110", "1111000000110011", "1110110101100100", "1110100111011111", "0000100110010110", "0001101101111100", "1111110110011101", "1111111010000100", "1110101111001111", "1111101011111001", "1111111000101011", "1111101110000111", "0001000110011010", "0010000000111001", "0000010110011001", "1100110110111110", "1111011000001000", "0001001100110010", "0001101001100100", "1110110111110110", "1110011101001000", "1111101001110100", "0000101110001100", "0001101111001001", "1111010101000000", "1110011000011110", "1110111100101001", "1111001100111000", "1111111111001000", "1101000011110111", "1101100001001111", "1100101100110101", "1111101111011011", "1110110110001001", "1111010101011010", "1111011110110010", "1101110111111000", "1111100001110001", "1111001011101000", "0000010010100111", "0001000110001101", "1111101100110100", "1111010000001110", "0000000011100010", "0000001010010111", "0001110101101101", "1111111011011001", "1110101000010111", "1110100011101001", "0000001011110111", "1110110001001001", "1111111001010100", "1111101111000001", "1111010100011000", "1110001110011001", "1101111110111011", "1110100001011011", "1111100011001110", "0000110000111001", "1111001010111011", "1110101001000101", "1110101111011100", "0000000000111011", "0000000011001000", "1111111100111100", "0001101011000001", "0000100000101101", "0001010100101011", "0010001101101000", "1111100010100101", "0000101100100011", "0001001011101000", "0001000101110111", "1111111011001000", "0001000001011100", "1111110110111101", "1111011000001000", "1111101111010001", "1110110010011000", "0001000101110101", "0000001111011001", "1111011011011010", "1110101111011100", "1111010111001000", "0000001100011100", "0000000011010111", "1110111001000000", "0000111010000101", "0001111001100100", "1111011101101011", "1110111110110110", "1111110011100111", "0001101111011100", "0001111011001001", "1110001011001011", "1111111011101000", "1110011011100100", "1111010010010010", "1110100100101010", "1110011010000011", "1101100001100100", "1111000111010101", "1111000010111010", "0000010101010110", "0000000101111000", "1111010001101000", "1110101101010101", "1110101101010001", "1111010000000100", "0000110011110100", "0001110110000011", "0010101011000100", "1110101110101111", "1111110001101011", "0001001101111101", "0000010000111110", "0001101000011110", "0000110111000101", "0001000001000111", "0000001101100010", "1110100001000001", "1110010001110101", "1110110010011110", "1110011100011111", "1111001011111101", "1111011101110011", "1110100011000010", "1110001100100101", "1111100000001010", "1110010100010100", "1111010011011001", "1110111100100101", "1111000011000001", "1110110011011011", "0000110011001010", "0000111101001101", "0001110100111101", "1111110001011000", "0000010110101001", "0001010000101001", "0000101111000010", "0001110100011100", "1111110100110110", "0001100010001001", "0000100101101110", "0000011001000011", "1111101011111100", "1111100111111011", "1110001010110011", "1111101101100000", "0000010101001101", "1111011000010001", "1101111010010100", "1111010001010100", "1110100111011110", "1110000101111110", "0000110101011010", "1111110000000011", "1111111101111110", "1111100110011110", "0001000101110111", "0001101111001110", "1111100110010101", "1111101010100001", "1111011111100010", "1111011100101110", "0000000100010111", "0001111100101110", "0001000110100111", "1111111010010011", "1110110110110101", "0000111001000110", "0000100101011100", "1111010011000100", "0000011001001001", "1111101000000100", "1110011111111111", "1110101010110100", "1111100110000000", "1111010100100111", "0000001101101111", "1111010011101110", "1110100000100010", "0000000011110001", "1110111010001100", "1110000100100011", "1101110010111100", "1111001001101111", "1111111111100110", "1111011000011000", "0000111001101001", "0000110010001110", "1111101011101110", "0001000001100100", "0000101100110011", "0010001010011101", "0001100111110001", "0001101010010000", "0000010100011000", "1110110011100101", "1111010000000110", "1111001000110010", "1110011100010100", "1101110101010111", "1110101111110010", "1111110010011000", "0000110001101011", "1111111011100100", "1111111000010010", "1110100100000010", "1111100010000000", "1111010111100000", "1110001111000001", "0000110111000101", "1011111011011110", "1101100001010101", "1110110111000110", "0000000111001000", "1111101110111110", "1111100000101100", "1110001011010010", "1110101001100010", "1111000011111010", "1111010001011011", "0000100001010000", "1110000111011000", "1111110111011100", "0000001110111101", "0001101011010110", "1110101000010010", "0010100000101101", "0001110001101101", "1110000110011101", "1110101000100101", "1110010000011001", "0001100101101000", "0001010110011111", "0000011111100001", "1111101010000110", "1101110110100110", "0000100001111100", "0010010101011101", "0000010011001110", "0001010101101011", "1101011010001101", "1101111011011110", "1111011010110101", "1110011011111110", "0000100100010001", "0000001001110101", "1111011010101001", "1111100011110101", "1111110010011111", "1110011111110000", "0000101111100100", "1111111001111101", "1110100001101011", "1111110000011101", "1111010110100000", "0000111100100100", "0000010001011000", "1110110010011001", "1111000000001101", "0010111000010000", "0010011011100100", "0001010001110011", "0000111100000111", "0001011001000000", "0001101111001110", "1111110011011010", "1111100101011101", "1111110101101110", "0000110110011111", "1111000100111001", "0000110100011111", "1111011111011111", "1111000100010111", "1110111011101001", "1111011010110010", "0000101000000001", "0000001010000100", "0000110110010111", "0000101010010101", "0001001111000010", "1101101000111100", "1110011101101001", "1111011010100110", "0000011000011110", "0001100111010101", "1110001110100110", "1101101101101011", "1100110110001110", "1110111101111010", "1111011100111011", "0010000010001011", "0000110001111000", "1111100010000100", "1110111001101101", "1101111110100000", "0010000111110110", "0000010111001111", "0000011111110111", "0001011011111011", "0001011001101110", "0000101101010100", "0000001011110101", "1111011000100101", "0000100111111110", "1111101000001011", "1111010100111000", "1111011110111011", "1110111111101111", "1111010100111110", "0000000111010001", "0000010010001000", "1110101011101110", "1110000010110000", "1101000010111000", "1110100011100110", "0001000111010111", "0000110100101100", "1111001100110101", "1110110000011110", "1100110010011101", "0000101001000001", "0000111011100101", "0000011000111111", "0001101001111100", "0000110101100111", "1111111101101000", "0000000001111011", "1110011111010101", "0000101110110111", "1111010010100110", "1111101000001111", "1110101101001101", "1111101100010110", "1111100111000111", "1111100101011100", "0000100001101111", "0000001011001111", "1110111110101100", "1110011100110111", "1101110101101110", "0000110000010100", "0001110100011000", "0000110000110100", "1111101011001010", "1110000110001100", "1110111000010011", "0000010100100001", "0001101101111110", "0000100011100010", "0010011011111111", "1111011101011010", "1111100001000111", "1111111000111010", "0001110010010100", "0000111101101010", "1111100000000000", "1111011000001101", "0000000010001111", "1111011110001100", "1101100101111110", "1110111000111110", "1110001110111010", "1110101101011010", "1101110100101010", "1101101110100111", "1110010001100111", "1111011010010000", "1110011011101100", "1101110100000111", "1101111001100110", "1110100000101000", "0001110011011011", "0000001010110110", "0000000000011010", "0000000101101110", "0000100001101100", "1111101110110001", "1110010110010010", "1110010110101111", "1110010101110010", "1111110101110111", "0000011001110111", "0000000010011010", "1111100110010000", "0001111000111100", "1111011111000001", "0000011011011000", "0010001001101111", "0010110000111101", "0001101000101100", "1100101011010001", "1110000001111111", "1111001010100001", "1111101001000100", "0000001101110010", "0000101100100101", "1110001101000111", "1110001010110001", "0000000011010101", "1111110110110000", "0010101100001110", "0000011010011001", "1111001011100110", "1111100010011010", "1110101101111101", "1111111011000011", "1110010100111001", "0000101100101110", "1111001101011100", "1110111010000111", "1111100101111110", "1110101110010111", "0000101001100110", "0000011101111111", "1111100011000011", "1111111010000101", "1110111111101001", "0001001110101011", "1111101101111001", "1111110101100010", "1110101011001011", "1101010110100100", "1110001101001101", "0000001001010100", "1110001011010100", "0000100011100000", "0000111111111000", "0000111111100101", "1111100110010100", "0000000000101111", "0000110001111100", "0010000101111000", "0000010101101111", "1111010001000010", "0010001000001101", "0000000110001010", "0000100000100000", "0010010101010111", "1110010100100101", "1111010110100011", "1110110010011101", "0000001000101010", "0000001101011100", "1101101100101100", "1110110000010101", "1111000100101011", "1110101011000011", "1111100111001000", "1111010001001011", "1101010000101100", "1111010101110010", "1110110101000011", "0000011111100101", "1111011111000111", "0000110101111011", "0000010000101100", "1111101011011101", "1111101010100101", "1110110101000011", "0000010111110011", "1110011101111010", "1111001110001111", "1111110010010100", "1111111011100011", "1110100010000101", "0000010000101000", "0000011100000110", "0000011100111011", "0000101110010101", "1111011010101110", "0000010100110111", "0000001001000100", "0000001011110111", "0000101011101110", "0000100101100001", "0000100101110100", "0001100100110000", "0001000100000010", "1111010110011111", "1111010000111000", "1111110101001010", "0000100001010000", "0000001000100001", "1110011001101001", "1100110111010011", "0000011011010101", "0001001011111100", "1111110111110110", "1111101000000010", "1110011111111011", "1111101100001010", "1111001110110100", "1110000100011010", "1111000111100001", "1111000000000110", "1110011100100110", "1110010011111010", "1111010010010000", "1111000110100101", "1110011010110000", "1111000101100101", "1111100001100000", "0000110010100010", "1111111110011101", "0000110000100011", "1101110010100111", "1101110010100100", "0000110110111111", "0001010101011101", "1110110000011111", "1111001100100100", "1111100011001000", "1110101001010010", "0000111000101000", "1110111110001000", "1110001011011101", "1111001110101101", "1111001011110101", "1111001011100001", "1111010001011010", "1111001101011011", "1110111111001011", "1111011100000110", "1111101110110100", "1110010111100101", "1110111000101100", "1110001100111011", "1111010101001110", "0000001100001101", "0001010010010111", "1110101111001011", "1110000110111110", "1110100000011110", "0000101010011101", "0000000011111100", "1110011110110010", "1111101101001010", "1110110111001110", "1111101000100001", "0000010010111010", "1101101111001001", "1110101011010001", "1110100001000010", "1110001010001110", "1111101001001100", "1110010101111011", "1111100000001000", "1111110010011001", "1111010001100001", "1111110110111101", "1110010010100011", "1110101001000000", "1111100110001001", "0001010010001110", "1111001010011001", "1110100001101001", "1111010110001010", "0000001100010110", "0010100001111010", "1111110101011101", "1111101101000010", "1111110111111000", "0000100011101101", "0011010000111010", "0001100010011010", "1110110010001001", "1111010110110001", "0001100001001111", "0010000010110110", "0000000010111001", "1111011111011101", "1111110011111110", "0000001110100110", "1111001000101110", "1111010111111000", "0000000011100010", "1111110000101011", "0001101000010000", "0000110100110000", "0000011111011010", "1111001001110010", "0000100111010001", "0000000000100010", "0001100010011010", "0000011101111010", "1110010100111011", "1111000111010100", "0001001101101001", "1111101101000000", "1111100100010001", "1111100011001100", "0001010110100111", "0001011000100001", "1111011011001110", "1110110000101111", "0000110001110100", "1111010011110110", "0000010011010101", "1111000001110101", "1110100101101100", "1111101100110110", "1111000001111110", "1111011110101100", "1111111010000101", "1110100000110010", "0001011001111000", "0001110100110001", "0000111001100110", "0000101010110000", "1111000010010011", "0001010111111110", "0001101101010100", "0000011100000001", "0010000011010101", "1111101000111001", "1111011000101110", "1111110000111100", "0011000011000010", "0000111100000011", "0000001000000110", "1110100100001110", "1111110111000000", "0000110101110000", "0000000011100111", "1111100001010110", "1111111101101110", "1110111000000111", "1111011101110100", "1110011100011011", "1111100111011110", "0000000111001101", "1111100100110100", "0000110001111001", "0001011101010111", "0010001011011101", "0001001011111010", "1111001000001110", "1111111100110111", "0000000111011100", "0000001110111100", "1111101010010011", "1110110101011010", "1101111000010001", "1110011000010010", "1110001001010100", "0001100010000001", "0001000100010111", "1110110010001010", "1110001111001101", "1101101001101100", "1111011011000011", "1111100101001101", "0000100100000101", "0001010101100011", "0001010011011101", "1111101000110011", "1110101011010110", "1110101111011010", "1111010011110111", "1111111011100001", "1111011110100100", "1111000100000011", "1101101100000000", "1110110111001000", "1111011100001101", "1111011010011100", "0000011000000100", "0000100100001100", "0000000101111101", "0000000000110010", "0010001001001011", "0011010100010110", "0010101001111011", "0000011011001011", "1111010001010010", "1111010001011001", "1111010110110010", "1111011000010011", "1110110010000110", "1111011100011101", "1110101110001111", "0000001001000000", "0000001000100101", "1111001010101000", "1110110010110011", "1110111010101011", "1111111000111110", "1111110010000100", "0000111110001111", "1110011010100001", "1111110010101011", "0000001101001000", "1111100001110010", "0000000001110011", "1111001111101100", "1110111101000110", "1110000111001100", "1111001000110010", "1101110110111101", "1111011100001100", "0000001101111001", "0010010110000111", "0001111100000100", "0000111010000110", "0000110000101100", "1111111101101100", "0000100011011000", "0000001111001000", "1111101111001001", "1111010101001011", "1111101100000000", "0000010010100001", "1111100001001111", "0000101011111111", "1111011100101001", "0000010011010110", "0000111001111010", "1111111101101011", "1111100101011100", "1111011110001111", "1111101100010010", "1111110110111000", "1110010001000111", "1101111000011110", "1110001000000111", "1111101110010101", "0000110010000111", "0001011101101001", "0001010010000011", "0001111101100110", "0000010110011010", "0001100101000010", "0000100101101101", "0001110010110010", "1111100001010010", "1111110111010001", "1111001110011101", "1111001111000111", "0000000011000101", "1110111111101101", "0000110001100011", "0001010010001101", "1111001111011000", "1101111000010111", "1110010111100100", "0000000111000010", "0000010011100010", "1111010000000010", "1110101111100000", "1111011011011101", "1111001001001101", "1111101110111001", "0000010011000000", "1111010001110011", "1111010100110111", "1110111111100101", "1110110010101000", "0000000011100100", "0000011010101011", "0000001010101011", "0000111001100011", "1111001010111011", "0000010011001001", "0000100001110100", "0000001101111011", "0000000111000100", "1111000111001110", "1110001001100001", "0000010111011110", "0000101010001000", "1110001100100101", "1111001011100000", "1111001000001110", "1111001101111010", "1111110000010010", "0001100000110100", "0000010110101110", "1111110110010110", "1110111010101111", "1110101000011000", "0001011100100000", "0000110111010101", "1111110111110101", "1110111010010100", "1110010000011101", "1111000011010011", "1111010001111111", "1110111110011110", "1111100001010010", "1111010000010110", "1110101011100110", "1111011100101001", "0000011100110111", "0000101010001000", "1110111111000100", "0000100111011111", "0010100111001110", "0001010001100001", "1111101011010011", "1110111111100100", "0010000110001110", "0010100011111101", "0000111011110111", "0010010111101111", "0011010010110101", "1111011111010011", "0000110001010011", "1111001011110100", "1111011010111111", "0000001001000110", "1111000001100001", "0000100011001111", "1101011011000010", "1100011010111100", "1110010011011000", "1111101001100100", "1110010110110000", "1110011000111010", "1110001100001000", "1101011001100110", "1111101000010010", "1110110001100001", "1110100101000100", "1111010010011100", "1101011001000001", "0000110110001110", "0010010110000110", "0000101111001101", "1111001001000000", "1111000100001101", "0000111001010001", "0001010010001111", "0001100001110101", "1111110111010101", "1111010001011111", "0000000100011100", "1111010010111100", "0001110001001101", "0010100010110101", "1110111001000010", "0000011110111101", "0000000101001001", "0000011100110011", "0001110010100000", "0000010100111100", "1111111101111100", "0000000000011001", "0010001111011110", "0000001111010001", "1111101110100110", "1110010110110011", "1110010001011010", "1100101101001101", "1110011010111001", "1110010001001110", "1110111100111111", "1110001110000010", "1101111110100101", "1111011101101011", "1110111110000011", "0000001110010111", "0000100010010001", "1111110101011010", "1111010100001001", "0001010101000100", "0001000101100000", "0000011010101000", "1110110010101001", "1110100110000111", "0001101000100100", "1111100011100010", "1110110000100100", "1101111110101100", "0000010110110101", "0001010100101010", "0010011111100101", "0000000101110101", "0000011110110010", "1110110010010010", "0000001110000000", "1111101000010111", "1111001101001001", "0000101110010011", "1111000001010101", "1111100011001010", "1111001101011100", "1111110001100111", "1111001110010100", "1111111100010101", "1110100011111010", "1111011111001111", "1111110010000110", "1101110101010011", "1110100011110001", "1101000001111011", "0000000111110111", "1110001111100000", "1111110110110010", "1110110001010100", "1110101010110000", "1110111110001001", "1101110101011101", "1111101011000000", "0001010001001100", "0000111001010110", "0000101001001111", "1110011011010000", "1101001010000001", "0001000101111000", "0001101111101011", "0000001111011101", "1111111010001011", "1110001011100010", "1111110111111100", "0001010110101000", "0001001110101100", "0000100000001110", "1110101111111010", "0000000110100000", "0000010001111100", "1111110010110011", "1111110011101010", "1111111010001101", "0000010100101111", "0000000011111111", "0000110110011101", "1110101010100100", "1101010000001001", "1111010111010100", "1111011101111110", "1111111100111111", "1110101010111100", "1101000001001000", "1110010000010000", "0000111110100000", "0000100100101010", "1111000100010001", "1101111010100110", "1111000110111100", "0010101011111000", "0000110000110000", "0000101111100011", "1111111111010100", "0000010111100110", "0000110111100111", "1111011100110100", "0000100100100001", "0000010011111110", "1111110111110011", "1111101011111011", "1110110000101101", "0000111111111010", "0001101011010011", "1111111011101110", "0000001000010100", "0001000011111110", "0000100010010001", "1110110110111101", "0000011000101000", "0001010001011011", "0001010101101010", "1111000011101110", "1110110111110010", "1111011100101001", "0000111111001000", "1111001100101001", "1111101111000110", "1111011011011111", "1111100101110110", "1110010001110101", "1110101111010001", "0000111011111100", "0000000000000101", "0001001011011011", "1111111000100111", "0000100111011100", "1111111011110100", "1111001111010011", "1111110101010001", "0000111111001111", "0001000010101011", "0000100111100101", "0000101101100011", "0000011011100101", "0000011001010100", "1111100101100111", "0000010100100101", "0000011110110100", "0000101001000001", "0001100110010111", "0001011110011111", "1111011111100110", "1111111000010000", "0000110010101011", "0001100111100011", "1111001111010010", "1110101110000000", "1110001001111011", "1111011101001001", "1111011001000011", "0000100110111101", "0000010110010111", "1111100001001101", "1110010001011011", "1110110001011101", "0000011001011001", "0000000111000011", "1110111001000110", "0001000000001101", "0000101110110110", "1111010100101001", "1111011001101001", "0000001011111010", "0010010010111001", "0010010100011111", "1111001101100011", "1111001101001110", "0001100010101001", "1111111000001000", "0000100011001110", "1110100100111001", "0000000111001010", "1111111011001111", "1100110001001010", "1101000101111001", "0000001100100100", "1111000100000110", "1110011011001110", "1110000011101101", "1101101001000000", "1111001111001000", "1101100111000001", "1110010100111011", "1111011110111101", "1111010000001000", "1110111101001000", "1111011000011111", "1111111000000100", "1110111011110100", "0000110011011111", "1110100001101100", "0000111011110011", "0001000111000111", "1110111100111011", "0000001010101001", "0000000110000111", "0000001000100011", "1111000000111001", "1110100111010000", "0000110110101101", "1110010110011001", "1111111110101101", "1111010110111100", "1111110111110111", "0001101111101000", "1110011010101011", "1110101010010100", "1111011111001110", "1110111110111010", "0001000011101011", "1110110011011010", "1111001001110010", "1111011110011100", "0000110001001100", "0011100001010000", "1111000100111001", "1110011110000010", "1110101011010001", "1110111101011011", "1111100001101010", "1110010110111100", "1101100110001100", "1110111000000100", "0000000110100101", "0001010010110011", "0000011100111011", "1110010001010110", "1110110110111101", "1111100111001110", "0000100001010001", "1111110011010011", "1110010100101110", "1110111100000001", "0001101010100111", "0010011000101010", "1100110101010110", "0000000000101000", "0001010010001111", "0001001100011001", "1110100111111110", "1110001101001111", "1111000001010101", "0000001111101111", "1111010100010001", "1110000101000011", "1110010101111011", "1111000110001101", "1111011000001100", "1100000100011111", "1101111010100010", "0000110000000111", "1111100001000110", "1110100111111110", "1111001111011101", "0001111000101010", "0000001111010011", "1110111011100010", "1111000100001110", "0000100000100111", "0001100011010001", "0000001001010101", "1111000110011010", "1111010001111010", "1111111110000110", "1111101010110000", "0000001110001010", "1111011101101011", "1111001000101011", "0000100101010001", "0000000000001100", "0001000110010111", "1111010111001100", "0000011001101101", "1111011001110101", "0000010010100101", "0000100010011100", "0000001010000010", "1111111100011010", "1111111110110000", "0001001011000011", "1111010001110111", "1111110111001101", "1111111110011111", "0000010100110100", "0001000100001110", "1110011101011000", "0000010011101110", "0000100110111001", "1111101100000101", "0001101000010001", "1111100100000100", "1110111100000001", "1110101000100101", "0000101010100010", "0000010010011001", "0001000011100011", "0000011100111111", "1110110100010001", "1111100101101011", "0000001100110000", "0000110000101000", "0000101100111010", "1110100001100011", "1101011000010110", "1110100111110010", "0001111111110111", "0000111000111111", "1111000001011010", "1101110111100000", "1111100011100010", "0010101101010001", "1111111010100000", "1110111010100111", "1111110100000100", "1110101110110100", "0001000100000011", "1110101010101110", "0000010010110000", "0010111010000000", "1111111101010011", "1111010010010001", "1110101010000101", "0011010100101110", "0000101011000001", "1111111101001101", "1110100111100011", "1110100101000010", "1101111101110011", "1110011101110010", "1110010001111110", "0000001111100011", "1101100010110111", "1110110100100000", "1110101100011110", "1111110100011010", "1110101110101001", "1101001111011000", "0000001000011111", "0010000010110011", "0011010110110100", "1110100101100000", "1110101100100101", "0001001100100001", "0000011001110101", "0000010101101110", "1101011000111011", "1111110101111000", "0000101100001100", "0000000101110001", "1111101001110010", "0000001101010110", "0000101111001110", "1111111011101011", "1111110100010010", "1111001000000000", "0000011000011100", "0000101100001100", "1111010011011110", "1111001011000001", "1110000110100110", "0000000111110010", "0010011011110101", "0000010000111111", "1110101010001000", "0000110111001111", "0001001001001010", "0001010001000100", "1111001011111111", "0001110011100011", "0000100111000101", "0000010010001010", "1111111011011010", "0001111101011000", "0000010110010100", "0001000011111100", "1111000100011010", "0000011000000010", "1110111111101100", "1110111101001110", "0010000100100110", "0001001010111000", "0000000111001001", "1110100011011011", "1111000001001101", "0001101110111100", "0001000010110010", "1110000001000100", "1111011000010011", "0000110110001010", "0010110000110100", "0001001101111110", "1110100011101010", "0000100111000011", "1111101011010010", "0010100001100101", "1110000111010111", "1111001101011100", "1111110101011000", "0001000001111000", "0000000011111111", "1111100011100000", "1111101011001011", "0000001001010001", "0000100110111011", "1111101101000001", "1110011100110011", "1101110011110000", "0000011110000001", "0000000010100010", "1111001110010000", "1110011011010100", "1111011000100110", "0000011100010111", "1111101101011000", "1101111100110000", "0001001001000100", "0000100010111101", "1111101110011010", "1110010001100001", "1110011001011000", "0001011001001111", "1111111010111101", "1110100111011001", "0000001000000111", "1111101110001100", "0000100101100001", "0001001011111001", "0001110011100000", "0000110000000010", "0000001100101110", "0000001101011010", "0000011000000011", "0000000101101001", "1111000101111010", "0001000010100111", "0000001111001000", "0000101001110101", "1110100101110001", "1101111101001010", "0000110011010001", "1111000110001110", "1110001011011010", "1101111100101010", "0001100101000000", "0010011000000111", "1110111010110001", "1110101000110101", "1110100001010101", "0000011110010101", "0000101010010111", "1111000001011010", "0000111100000000", "0001111101000001", "0010101101110101", "1111111010110111", "1110010110101011", "1111000111110000", "1111110111110100", "1111010011110101", "1110001111111101", "1111111111011001", "1111001110011001", "1101101101100011", "1101111110101111", "1101101000111100", "1110011010001111", "1110000001011101", "1101111011000101", "1111001001110000", "1110110010010010", "1110111100000101", "1101001110000001", "1101001011001010", "1111110010001110", "1111101000111000", "0001000100111111", "0000100001100010", "0000111100000100", "0001011110010010", "0001101000101101", "1110110000010110", "1110111001010100", "1111101000010011", "0000100000101000", "0000011001010001", "1110100011011011", "1111100001000000", "1110001010101110", "1111000111001000", "1101110101100101", "1111010101011000", "1110100100100110", "1101110011001010", "1110100111000011", "1111100010100011", "1101111101001000", "1101001111101001", "1101010101111110", "1110111100001110", "1110110010110101", "1111101000100010", "1110100011101110", "1111110110000000", "0000101111100000", "0000001001111001", "1110010100000100", "0000001011101101", "1111101110110110", "1110111000011001", "1111011100011001", "1110100110010000", "0001000010000010", "0000110000101110", "1111111110101010", "1110111000101111", "1111001110001011", "0001001100011000", "0000100111111100", "1111011111011010", "1111101111111010", "1110011001011001", "0000011111110111", "1110110001010001", "0001000111101010", "0000010010010100", "1101101110111010", "0000101000001101", "0000010000110011", "0000001001100111", "1111000000110111", "1111011001111110", "0001010101010100", "0001011010110100", "0001001101000010", "1110100100010110", "0000100101100011", "0001001000101110", "1111111010111010", "1110010010101010", "1111100110111100", "0001100000110101", "1111111111110000", "1110000011101011", "1110110101011100", "1111101110111110", "0000110110001010", "1101011110011111", "1110110010101100", "0000000001101001", "0001001011110100", "1110001101010000", "1111011111101000", "1110010011001001", "0000010101110010", "0000101110101110", "1110101001111000", "1111111100011001", "1101100110000111", "1110000110110101", "1110011111010101", "1111100000011000", "0000100001010111", "1101100000100101", "1110101010011010", "1110001101010010", "1111001111111000", "1111001111101010", "0001101001111111", "0100010000101110", "0000110100101100", "1111111011100100", "0001110001111100", "0011000101010110", "0000100000010111", "0000010111111111", "1110000101010111", "0001001100010100", "0000100001001000", "0001011110110000", "0000101100111010", "1111110111001100", "1111001001100101", "0001001010101001", "0010010011111101", "0000110111111111", "1111110010000110", "1111110101010000", "1111011101111001", "0001110111011101", "0001001101011111", "1110011111100100", "1111110111000110", "0000110110001110", "1101110101110000", "1111010110101101", "0000110110000011", "1111101001001100", "1101111010100000", "1110100010100111", "0000110111111100", "1110101101001111", "0000010110101011", "0000110011110111", "0000110001000010", "1111111001101010", "1111000111010001", "1111100000101110", "0000001001101110", "1111001110111000", "1101000001100011", "0000111101110001", "0001010000101011", "0001011111010011", "1110010110000110", "1110011001101101", "0001100111101111", "0000110110110001", "1110110101100100", "1101110101110010", "1110100010001101", "1111011001000101", "1111001011001000", "1101100110001111", "1110000011001100", "1110110001010000", "1110010001101010", "0000000100111101", "0000011000011101", "1111111011000111", "1110110100000010", "1110100110101101", "1111100101110010", "0000001110101011", "1111111011001010", "1110100110000001", "1111010001111100", "1111001101000101", "1111110101101110", "1111011111001110", "1111111110010010", "1110011110011110", "0000000011110001", "0000011010101000", "0001100000001110", "0011000000101000", "0001000011000101", "0001110110000100", "0010001100100100", "0001100010000010", "1111011000110001", "1111110101011101", "0000110100101110", "1111111100100101", "1111110010000111", "0010010011000011", "1111101101010000", "0001110011000000", "0001011101011000", "1110101110001001", "0000100001100001", "1111001010011100", "1110100000110000", "1111011010101000", "1111101010000110", "0000101010111010", "1101011010010101", "0000110001011000", "1110111101001111", "0000010101110111", "1110110111100111", "1111100011111011", "1111011101110001", "1111101001101011", "1111111010001000", "1111000111110101", "1111110101100010", "1111111111011001", "1111110011011000", "1111011001110000", "0010100000101011", "1111110010110101", "0001011000100011", "0001010110100100", "0000011011111001", "0001110111101001", "0000011010010100", "1111010110001101", "1111111101011111", "1111001010100100", "1111010001011010", "1110111101010000", "0000001100101000", "0000101111100001", "1111010010000111", "1110010000101111", "1111000011010101", "0000101010110011", "1110110110000000", "1101100110100110", "1111100001110101", "0001101010000011", "1111111011111110", "0001001111001010", "0000000100010010", "0000100100000001", "1111001001001001", "1111100111000100", "1111110111101011", "0000111010110011", "0000011000000111", "1111010011010101", "1110000001011110", "1101011110111111", "1110010011000011", "1111110111011101", "1100101010001111", "1101010110000000", "1100001101111101", "1100011111000000", "1101101011011001", "1101001111110110", "1101000011110001", "1101011010100111", "1111001011011011", "0000111100010000", "1110011010011010", "1111010001101010", "1111111000101110", "1111010110010111", "1111101101110101", "1111001111001110", "1111100011001101", "0000101100010010", "1110110111111111", "1111001010111110", "0001001101101011", "0001010011000011", "1111001011001101", "1111010011111101", "1110011010100000", "1111110011010111", "1111011110010001", "0000011001101001", "0000110100110000", "0001001111100110", "1110011110011001", "1111001011000011", "0001001011010100", "0000110010101111", "0000001101010101", "1110000101111000", "1111110100101111", "1101110001100101", "1110110010110110", "0001010011101101", "0000101110010000", "0000011100001000", "1110010011001101", "0000010110011110", "0001101111101101", "0001000111111011", "0000000001100000", "1111001001111011", "0001000010001001", "0000000101101001", "0001111010111101", "1101010101110111", "1111010001111010", "1110110101001010", "1110010000011010", "0000001001011010", "1111001100111000", "1101000100011011", "1100101010010110", "1111000100011011", "1111110101010011", "0000111100110100", "0001011001110110", "0000010100000010", "1110100011011101", "0000000011000110", "1111011111101101", "0000111100101000", "0011010011011100", "1111001000001001", "0000110100101101", "1110101111000011", "0001001000101101", "0010011000100110", "0000001011100010", "1110110001111111", "1111111101100000", "0001000010101000", "0011100110110111", "0000100100111111", "1110111101010001", "1110111011010000", "0000000001110001", "0001101010001000", "0000000100101011", "0000110100000001", "1111110110111010", "1111001011011000", "1111011110001011", "1111010011101011", "0000111110011111", "0001100010110010", "1111110010110000", "1111110110100101", "1110100101101010", "1111010100111111", "1111110000111011", "1110011100011001", "1111000000101110", "1101000110001110", "1111000101010100", "1111001011101011", "1111010000100000", "0001001100100101", "1110110001111001", "1110001011110110", "1110110100111100", "1110110011011101", "0000110011000111", "0000001001010101", "0001111000010011", "0000110111010011", "1111101110011101", "1111100101010101", "1111011100100111", "0001000101011111", "0001010100010101", "1110011100110010", "0000111100011010", "1111010011000011", "0000010111111011", "1110110000110010", "1111000010000111", "0000001010000111", "1110101011101101", "0000010000011001", "1101101101011110", "1101111100111110", "0000001010011011", "1111000101010000", "1111100101100010", "1110010101010111", "1111100110011010", "1111011101101101", "1101111001110010", "0000010100100100", "1110100100011111", "1111001111000000", "1111001110010010", "1111011110110100", "0000011010000000", "0000101001011001", "1110110111101100", "1110110100011001", "0000110110010011", "1111000100100010", "1111001111010100", "1101110101011111", "1111110001000001", "0001011000000100", "1111010010010001", "1111000100010001", "1110110100110010", "1111111000000110", "0010111110110110", "1111001001101100", "1111011010100101", "1111111001000101", "0000001100001101", "0001000111010001", "0000101101100110", "1111111110010101", "1101100001011010", "1110011000101010", "1110111111010110", "0000111010100110", "0000001111001010", "1111100100101111", "1101110001111101", "1111100110111101", "1111010010111110", "1111001010000111", "1111011010100011", "1110010100101100", "1110110011001100", "0000000101111111", "1110111100011010", "1110111000001001", "1110111000000010", "0000111011010011", "1111110000011110", "1110100011101010", "1111001011101111", "0000100000111010", "0001011111000110", "1110010111110111", "1110001110000001", "1101001011001010", "1110100101011100", "0001111101000010", "1111001110010010", "1111111001001001", "1111100101010001", "1111011111101000", "0010010101010000", "1111101100100001", "0001010001100011", "0000000101010100", "0000100100000001", "0010100100001011", "0000110100010000", "0010010100110110", "0001001010110001", "0001010001100011", "0010111011111100", "0001100000010011", "0000100100000010", "0000110001111011", "1111010100111001", "0000001001000111", "0000110000101001", "1111100011100000", "0000101110100111", "0000010001000101", "0000010110011011", "1111100111100110", "0001101111000001", "1111111000001010", "1110110110011000", "0000001001100100", "0000111110001000", "0000010110010010", "1111111101111100", "1111111110000000", "1110100000000001", "0000100111001000", "1110010000010111", "1111000000001111", "0001011001101110", "1110100011111101", "1111101111010100", "1101011010010011", "1110010011010111", "1110101010111010", "0000000010000110", "0000011111000100", "0000101000000010", "1111101101001000", "1111111000110001", "1111001000101111", "0000110111000110", "0001001100111110", "1110101110101001", "1111001110111101", "1111011100001001", "1111100111000000", "1110111110111101", "0000001100101000", "0000001101111011", "1111110000100011", "1110010100001100", "0000001101100010", "0001000100111001", "0000111011001100", "1111100111001000", "0000010011000110", "0010001001001001", "0000110100000100", "0001001111000011", "0010101010100010", "0000001001110000", "1111011100100111", "1111010010010011", "1110111001001101", "1111100110100011", "0000100010101011", "1110110010110110", "1111111101011001", "0000001000000111", "1111101001011110", "0000110101000110", "1110001001100011", "1111001110000001", "1111011001111111", "0000011110010101", "0001011100000111", "1111110101100011", "0000011010101011", "0000100111010000", "1111011001010000", "0000111110110100", "0000010111100010", "0000111001011100", "0001010100010100", "1111111110011001", "1111010100001011", "1110101000001111", "1110100011000100", "1110011001101000", "1111110001111010", "1111001010011111", "1110101111011011", "1111010111111001", "1111100100100000", "0000001001000000", "1111101000111101", "1111110010111110", "1111100000100101", "0000001010111001", "0000100001100111", "1110111110011100", "0000100111100010", "0001010100101101", "0000010010100111", "1110001010001011", "0001001000101010", "0001110100110101", "0010100011001011", "1110100000001110", "1100110111110000", "1111111111110111", "1111100110011000", "1111000101001110", "1111000001110001", "0000111111011110", "0000000010011101", "1111101011110000", "1111101010001001", "0000100100000011", "1111111010011010", "0000011101111001", "1111110011101001", "0000101100110001", "0000001110111000", "0000101111111100", "1111010110010001", "0000001100011001", "1111100100100011", "1111011011110000", "1111100001100111", "1110000100001111", "1110111001011011", "1101111110000111", "1111001010110111", "0000101110010110", "1111111100100000", "1110100000000001", "1110001110111010", "1111010001000001", "1111111110001001", "1110011001011111", "1110111101111011", "1111001111100011", "0000000001010011", "0000000100111010", "0000011001001000", "0010000101000111", "0000010000000011", "1111011101010110", "1111100010100111", "0001100001001111", "0000000110100010", "1110111011011010", "1110011001000010", "1111000111100111", "1110101110010110", "1111100110011000", "1110000001010000", "1110101100011010", "0000011110010001", "1111100111011111", "1111110110000100", "1110101001010010", "0000000010111001", "1111011001010010", "1110101001111100", "1111010010111000", "1110101011000000", "1111000111100010", "1111101100100111", "0001010110001000", "0001101100011111", "0000011101101000", "1111101110001101", "1111001011010110", "0000110110101101", "0000010111111111", "1111100111100000", "1110011110001001", "1111000011111011", "1110011110000010", "1110111101011010", "1110101101011000", "1101110011100110", "1111000101101001", "1111111110110101", "1111101110110010", "1111111010100111", "1110101101010101", "1111101110110001", "0000000110010011", "0000010000010100", "0000111001111001", "1111011001111011", "1111101101111111", "1111110001110101", "0001000110000000", "1111111101111110", "1111000010100110", "0000000001100111", "0000011001011000", "1111101110011111", "1111011111001001", "1111001101000001", "1111010111011101", "1111001100111001", "1111110100010110", "0000010000110100", "1111011000101011", "0000100000011001", "1111010000100110", "1110001000011001", "1110100101111110", "1111000001111001", "0000111100100000", "0000000000000011", "1110101001011010", "1110110110101100", "1111010010011100", "1111010000001011", "1111010001101010", "1111011001100100", "1111010110110111", "1111110011101101", "1111110001100011", "0000001001111100", "0001100001101101", "0001101000100101", "0000000000100101", "1111000100001001", "0001111000100110", "0001110001001010", "0000101100110110", "1101111110001100", "1111010111001100", "1110000101010101", "0001000111011111", "0001110101001011", "1110100101010010", "1111011111001011", "1110100111110100", "1111100111001010", "1110111111101001", "1111011000101111", "1111011101100001", "1111000001101101", "1111100001000011", "0000100110010110", "1111010101001011", "1110101101111111", "0000110001100011", "0000001101011001", "1111110001001100", "0000111001101000", "0000001010110100", "0001111000101110", "0001000110110000", "1110100111111000", "0010000011010011", "0001001100111101", "1110110001001010", "1111111101011000", "1111001010010011", "0000010000001101", "1110111110010110", "0000001000001110", "1111001100110001", "0000010100111010", "0000101011101110", "1101111110100111", "0000001001101001", "1111111110001000", "1111110101011010", "1111101100110000", "0000101101111011", "1111000010011111", "1111011101000001", "1111011001001000", "0000000011011010", "0000111111110101", "1111101111110110", "1101110001011011", "0000101101001111", "0000101111110000", "0000011010011100", "0001101000111000", "0010010010111000", "0000010101000100", "1110101001001100", "0000001011010111", "1111101110010010", "0000100111110101", "0000001111011000", "1111000011110001", "1110111101011101", "0000010001111111", "0000011111110100", "0001000000011110", "1111001010111011", "1110000110001110", "0000000100001101", "0000011110100100", "0001100100100111", "0000000111101000", "1111100101101010", "0000000100001111", "0000001100010010", "1110110001011100", "1110001011100110", "1110100110100101", "1111010011011100", "1111010110000011", "0000001100110111", "1110011010000111", "1101100000111100", "1101111001101001", "1110010101011001", "1110111111001110", "1111110011111101", "1110110000001110", "1110110100101001", "1111001011100101", "0000110100000111", "0000010100011001", "0001010100011111", "1111100011101100", "1111101011110110", "0000111000110111", "0000011101111011", "0011001010001011", "0000010010101000", "0000001101000010", "0001000011001010", "0011010001110001", "0011110000111001", "1111111100001011", "0000001101111100", "0000001100011001", "1111110010010100", "1110111110110001", "0000000011011101", "0000110000111010", "0000011111000111", "1111010011010011", "0000001110010100", "1111001000001111", "0000101001010101", "0000000110110111", "0000010011010101", "0001111110000000", "10000000000000000", "1111010100110010", "1111100100110001", "1111100000001101", "0000101110100011", "0000000100110001", "0000010101101100", "1110101101110011", "1111111010101000", "1111100101001111", "0001011000110101", "0000011001101011", "1111001100011111", "1111111001101000", "0000011001001001", "1110110000100100", "0000011100011011", "0000110010010111", "1110111100011100", "0000001101011000", "0000001010100000", "0000100101101111", "0000111111000011", "1111101011001001", "0000111111000010", "0000001001000010", "1111001111111100", "0000010110000000", "0000010011010011", "1111001001011100", "1111111000011111", "0000001110101010", "1111111111011001", "1110111010001110", "1101000010011001", "0001000111101010", "1111011011011010", "0001100010000111", "0001101100001011", "1111111100001101", "0000101100110010", "0000010001111110", "0000001000110000", "0000000111010001", "0000010101000010", "1111100001101011", "1111111001000101", "1111001101000000", "1110111011000101", "1111100100100111", "0000011010111110", "1110111001110100", "1111000001100111", "1110111110111100", "1110111111000010", "0000110111101110", "0000101110011011", "1111100010000000", "1111011001100111", "1111001010101100", "0001101100100000", "0001101100011001", "0000100011001010", "1101111101111010", "1110101101100011", "0000001000110100", "0000010101111111", "0000110111011011", "1110101100100111", "1110000000010011", "0000000000101001", "1111010001000010", "1111011011101010", "1111001100001000", "1110010011001001", "0000011101011010", "0000000111000111", "1111111111100110", "1110111100100110", "1110010001001100", "0000001101101001", "1111101011100101", "1110010100110010", "1111000001001000", "0000001101000000", "0000010011011010", "0000111100001011", "1111000010100101", "1110101000111100", "1111001110001001", "0001101000011111", "0001100000111101", "1111101010101110", "0000010111111110", "1111100011111101", "1111011001100000", "1111010111010000", "1111001000011010", "1110111101001101", "1111110110001111", "1110010101010001", "1110111111011111", "1111100101011110", "1110111011011001", "1101111100111100", "1111100111110001", "0000010011110100", "1110101101001100", "1110011111000011", "1110000110010100", "0000110000000000", "0000010000001100", "0001011000010000", "0001001101011101", "0000100010001011", "0000001000111000", "1110000000110010", "0000100011011000", "0000101010011101", "0001001010111000", "0001001100000000", "1110101000001001", "1111001111101011", "0000000001100110", "0000011000000110", "0000010011000011", "1111010010011001", "0000010000110000", "1110100111010001", "1111000000000001", "0000111101011110", "1111111011011010", "0000000010111101", "1110010110001011", "0000100100001010", "1111111101101010", "1111010100111001", "0000011000100001", "0000000110110010", "0000010101000111", "1111011000001111", "0000010110101110", "0000100111011110", "1111111101111111", "0000000101101110", "0001110110001100", "0000010010000010", "1110110110111111", "1111111100110111", "0000111000100111", "0001010001110100", "1111010011001101", "1110011010100000", "1111100110100110", "1111111111001111", "1111101100010101", "1111101011111001", "0000001001000001", "0000000001101010", "1110100000011110", "0010000100110011", "0000000011110110", "1110000110010100", "1110010110001001", "0000011001001101", "0000111010010101", "1110110011011111", "1101101101000000", "1110100001011000", "1111110010100010", "1110001100110110", "1110111000111000", "1110010110011011", "1110111000110100", "1111010111001010", "1110011110111000", "1110111011000101", "1110110101011111", "1111100011000101", "1110110100101100", "0000011000100011", "0000011101110011", "1111110101001110", "0000001000001110", "0001011111001111", "0000011011100001", "0000001000101001", "1111001000111010", "0000000001001101", "1110101010111000", "1111110001110100", "1111011011001010", "1110110101001000", "1110011010001010", "0000000101000011", "1111110000000011", "1111010100110011", "1111100010110110", "0000001111100100", "1110110100100100", "1111111000001100", "0000010110001111", "1111001101010001", "0000100010011010", "1110111001110010", "1111010111111100", "0000011111001011", "0000001111001011", "0000101001011001", "0001110000011010", "0000000011111111", "1110100101100010", "1111111011001010", "1111111001001010", "1111100010010000", "1110010000010001", "1111101001010100", "1111101110101000", "1110100101010010", "0000000010001000", "1111011111100010", "0000110000110010", "1111100001100000", "1111101010000100", "1111101111100001", "1111110111000010", "0000000110111110", "0000011000010011", "1111101001000110", "1110111011001110", "1111101010001000", "1111101111000010", "1111101010111101", "0000001111000001", "0001111011010010", "1110011000110100", "1111111101111100", "0001001110111010", "1110100100101101", "1111111110100000", "1111111000010110", "0001100011001100", "0000010001110100", "1111011110011110", "0000011010110001", "0010000000111010", "0001001111110010", "1111000110111110", "1111011100101011", "1110111110001001", "1111011101010110", "1110001110100010", "1111011001111011", "0000001111101000", "1110011000000010", "1110001110000011", "1111000100110111", "1111001000000101", "0001011011100110", "0001100011000010", "0000100101101110", "0001110011001110", "1111011110111011", "0000001101000001", "0000101001100001", "0010000100011011", "0001000101010000", "1111111011111011", "0000000110010001", "0000110011110111", "0001111000000111", "1111001110001101", "1101111001001001", "1111011010110111", "0000011111100011", "1111001111001011", "1110011111100001", "1111000100100111", "1110110010010100", "1111011000100100", "1111010010001010", "0000001001010010", "1111110011011101", "1111001100010101", "1110010100101011", "0000101111110001", "1111101100000110", "1110010101110100", "1110011011111011", "1110100101110000", "1111000011111110", "0001010010111101", "1110100100001011", "1110001110011100", "0000011101010011", "1111011011010101", "0000000011010100", "0001101000100000", "0100100001001000", "0001100110001010", "1110111100001111", "0010010100100101", "0010001001111011", "0010100000101010", "0000111011101011", "0000110101001111", "0000101000011011", "0010000101001110", "0001010010101011", "1111100110111011", "1111010001000011", "1111100011000111", "1111000000011001", "1101111001100101", "1110111000001000", "0000010001000001", "1111100000101101", "0000000101000011", "0001111001000101", "1110011010010100", "0000100010010101", "0000010000011011", "0010100101111111", "0001001101000001", "1111110110111111", "0001100110001110", "1110100110000100", "0001010000001101", "1111000100100010", "1110101000011111", "0000000001101111", "1111000101111010", "0000010000001001", "1110111011110011", "1110010100100101", "0000000100001011", "1111110110101000", "1111101101011100", "1110110100101000", "1110001101001010", "0000111110010000", "0000110000000110", "0000010011011101", "1111011011000110", "1101100100111100", "0000110000000010", "0001000010001101", "1111000010111111", "1110010111100010", "1111001100101101", "0000101010100101", "1101101010011110", "1101011001110011", "1110111001100100", "0000100111101000", "0000011101000011", "0000011000101011", "1110101010100010", "1110101001110101", "1101111100010110", "0000001011010001", "0000101110001011", "0000110001101001", "0000101110010000", "1110111101110101", "0000000010001010", "1111101101100000", "0000001000101001", "1110101000011101", "1110111110011101", "0000000001010000", "1110111110100000", "1101111000000111", "1110001011011111", "1111100110001101", "0000011000111010", "1111100110111011", "0001000100011010", "0000101001110110", "1111011011001001", "0000101111011101", "0000011011000110", "0000110100011100", "0000000101100011", "1111000100000001", "0000000110100011", "0001000100111101", "0000111011000111", "1110100010101000", "1111011001101100", "0001001001111111", "0000011000100011", "1111010011000010", "1110101101011101", "1111101101111000", "0000000011100000", "1110010111001010", "1111010100101110", "1111110011111011", "1111010000001000", "1111011100100011", "1110111000011011", "1111001010011111", "0000111011100100", "0000101011010010", "0000000111100110", "1110111011111110", "1111101010111100", "0001000100110110", "0000001101100100", "0000000101010110", "0000111110011001", "0000111110010100", "1111011101010110", "0000011000110010", "0000111010100110", "0000100101101100", "0000011001001101", "1111010101011101", "1111000101011001", "1111111001011111", "1111000001100001", "1111010010111011", "0001010100111100", "1110111111011011", "0001001110100100", "1111001011110111", "1101101110001000", "1110011011000010", "0001001010010011", "1111000100000111", "1110101110110110", "1110000111010001", "1110110110111000", "0000101010001101", "0000000011001011", "0000001111110111", "1110010100111010", "1110011100001001", "1111101101010101", "1110101111001111", "1110011010111000", "1101011011010110", "1110000110100000", "0000001111101000", "1101100000001001", "1101010101110110", "1101001001101000", "0000100101011110", "0001101000011001", "1110101001111100", "1110000001010000", "1110010001001000", "0010010100111100", "0011001100000111", "1111000001110001", "0000010110011000", "0010100111101100", "0010111001001100", "1101111110111001", "0000110110101101", "1111110010000000", "1110011011010010", "1110011000111101", "1101111101101110", "0000110001110010", "0001110110010101", "0000100100111001", "0000111111011011", "0000111100111010", "0001010000101000", "0000001111011100", "1111010010110110", "0001010111011011", "0001010001001111", "1110111111010000", "1110010101100101", "1111100110010101", "0000110101000100", "1110110111111010", "0001001010101001", "1111010111100101", "1111010000011110", "1111110000001001", "1111010011100010", "0001101100110011", "0000011110110000", "0000101000101110", "1111100111001110", "1111110001001110", "1111101100010000", "1111110011010110", "1111000101000000", "0000010100011010", "1111101111101010", "1110000110000010", "1111101110010011", "1111001110001111", "0000100010001110", "1111110111010100", "0000110011100010", "1111001010010001", "1110111000111100", "1110110111010000", "1101110010010010", "0010100000101000", "1111101010100110", "1110010010101011", "1111101010111011", "1110111101100100", "1111100001001100", "0000011000101000", "0000101101100100", "0000110110101100", "0001110111010000", "1110101100011011", "1110001001111110", "1110110000111101", "1111011000110111", "1111111101100111", "0000011100010000", "1111011001101101", "1111110011001011", "0001010110101000", "0000101010110001", "0001011011010001", "0000011011011111", "0000001111100000", "0001001001100001", "0000110010110100", "0010000111010101", "0000010001001101", "0000000100010100", "0010001110010101", "0001101111000010", "1111011001100000", "0001000100111110", "0000101000101100", "0001101011101101", "0001110000101001", "1111001101110001", "1111011111101101", "1111111010111011", "1110100011011111", "1110011011101110", "1110100001111100", "1111000111111001", "0000001001101111", "0001001000111110", "0001010101001000", "1111101101100100", "1111001011100111", "1111100001100110", "1111101001010011", "0000000010111101", "1111101111111101", "1110111000111101", "1110010100111000", "1101110100101111", "1110100010111101", "1111001110110000", "0000010101010001", "0000000000001000", "1111010001110000", "1111010010010100", "0000101011011010", "1111110100101000", "1111001110011101", "0000000011110000", "0000010101111110", "1110110111101110", "1110100100001111", "1110011111000011", "1111010111110001", "0000111110000111", "0000001011000110", "1111011000110010", "1101110000101111", "1111001110101011", "0001111100111000", "0001011101100110", "1111110110011001", "1101111111111000", "1111111000100011", "0000111100001011", "1101101001001010", "1111110110110100", "1111100111110100", "1110101011111101", "1111011101111001", "0000100101011000", "1111101000001100", "1111001000001101", "0000000010000010", "0000101011101010", "0000010101100011", "0001100000000100", "1110011001101001", "1110110011111110", "1111110011011011", "1110010100000111", "0000101101100100", "0000011011111011", "1111000111000101", "0001011010011101", "1111011001011000", "0000011000101111", "1110010010000101", "1111001101011110", "0001011110111010", "1110100001100000", "1111010101101101", "1111110010010110", "1111001000110100", "1111001100010001", "0000011011001001", "1110101111001000", "1111011111010010", "0000110010011111", "0000001111010011", "0000000000110001", "0010000101011101", "0000011100110001", "1110001000111101", "0000000010011110", "1110100110100001", "0001100100111110", "0000100010110110", "0000000000100001", "0000011111111010", "1111000000101100", "1110110110001100", "1110110011101010", "1110100001110011", "0001001010110110", "1110100000010100", "1110100110101111", "0000000010000111", "1110111000101010", "1111100100001111", "0000001011101101", "1111100100000010", "0000000101101001", "1111000000001101", "1111101011010011", "0001101101000010", "0000110010010100", "0000101010111111", "1111100000000000", "1111001010000110", "0000000000010111", "0010010100111001", "0000101111110110", "1111101000011001", "0000001010110001", "0000101000111100", "0010111111100011", "0000011010110001", "1110101001110100", "0000101001111000", "0000111010001110", "0001001110010100", "0001111000011011", "0001011111110010", "0001000110010010", "1111000100101101", "1110111111000011", "1110010001000011", "1110101100010111", "1110001010110000", "1110011110000111", "1111001101111101", "1111101010110000", "1111100101101001", "1111110001001000", "1111001101100000", "1111010001101000", "1110011010101001", "1111011110000111", "1111000101000000", "0000101001111100", "0000010011010110", "1110000011000110", "1110110000000010", "1111101101110010", "1101111000000101", "1111110010101100", "0000010001000001", "1110110101000111", "0000010011111101", "1101011101001001", "0001001000010111", "0001101111011001", "1111110100000011", "1110011010110001", "1110111101100000", "0001011000001110", "0001011000111101", "1111110010010110", "1111100001011011", "0001001101001110", "0001011010101011", "1111100011000110", "1110011100011011", "1111000110011000", "0000110100001110", "0000100000110101", "0000001011011101", "1111100111000110", "1111011101100111", "1110101101111001", "0010011001000000", "0000110000000111", "1111100101011100", "1110010110111111", "1111011101100000", "0011000000100001", "0000100100011000", "1111010001111011", "1111010010100101", "0000111000010011", "0010011111010001", "1111101011101000", "1110100111100010", "1111010010110110", "0000101010000100", "0001011010101001", "1111110110110111", "1101111010000001", "1111101011001110", "0001000111000110", "1111011111110010", "1110001000001111", "1110101010011010", "1111011110011111", "1111010101100110", "0000000110100110", "0000001111101101", "1110100011111100", "0000000111111110", "0000011001101001", "1111001000100100", "1110100010101010", "1111100110101111", "0000111101001010", "1110000010100100", "1110100101001111", "1101111100001100", "1110111111000000", "0000111000000001", "1110011011010100", "1110100010100000", "1111000001010010", "1111000001011111", "1110011110000100", "1101100011011000", "1111010001001010", "1111100010011110", "0000000100001010", "1111000010111110", "1101010111001101", "0000011000001011", "0000100000010110", "0000011010001011", "1110111011001001", "1111010101011100", "0000111101110011", "0000110100001101", "1110000101101011", "1111001101110010", "1111101111110110", "0010011011100010", "0000101000111000", "1110000101010000", "1110100100110111", "1111110110111100", "0010000001011110", "0000000000011111", "1101110000101100", "1111010101001000", "0010010110100101", "0000000111100101", "1111001001100110", "1110000110011011", "1111110111101100", "1101001101111011", "1100101010001111", "1111101110011101", "1111110000101000", "1110101101010011", "1101101111111110", "1110110100100000", "0000011111010100", "0000000011101100", "1110010011001001", "1111100101000000", "0000010000111001", "0000011010000111", "1111010010011011", "1111011000110101", "1110110110110000", "0000010110111010", "0000010100010010", "1110111110001010", "1111110110000111", "1111010010111011", "0000010000101001", "1111000110100110", "0000000111000011", "1110100001011010", "1110001010111101", "1101011110111001", "1101011101100110", "1111001101101110", "0000000110001001", "1111010011111011", "1110000000000101", "1111110010110100", "1110101111001001", "0000000101001110", "0000001000000010", "0000010110010001", "1111111000101001", "0000001101001111", "0001000111110010", "1110100110111111", "1111111011100010", "1111000110111010", "0000111010001011", "1111011101000001", "1101111110110010", "1111011110011000", "1111000110101111", "1111001100000011", "1110110110101101", "1111000010010101", "1110001011001101", "1110000100011001", "1111010011000111", "1110111011001011", "0000000011000010", "1101100010011101", "1111111001001100", "0000010000101110", "1111110011111010", "0000110001110010", "1110010111000101", "0000010101111001", "0001001001000101", "0000101111000000", "1110100000011000", "0001001011001001", "0001010101010000", "0001000011010111", "0000000101000011", "1110101101001011", "0010111010011000", "0001101000010000", "0000110000110001", "1111111110001110", "1110110100111010", "0000000011110110", "0000100001010001", "0000011110100011", "0000100011000110", "1101100010000100", "1110000000101101", "0000000111011101", "0001000011111111", "0001100100111101", "1100100010101001", "0000100011100001", "1111011110101010", "1110110111110010", "1111001111110001", "1111001011101111", "1111111100111110", "1111111111000111", "1110010101000011", "1111001111010100", "1110010101001110", "0000011010010111", "1110110111111101", "0000000110111111", "1111000101101100");
    Plus112_i_1 <= ("1111010101111001", "1111001000010001", "1110110111110011", "1110010111000111", "1110100100010011", "1110010001101101", "1110111011100000", "1110011011110011", "1101110110101010", "1101111011110011", "1111011001000001", "0000000110110011", "1111111101101111", "1100101011101010", "1110100100011110", "1111101100001110");
    Times212_i_1 <= ("0000101110111010", "0000111110001011", "0000101011101100", "0000111110110001", "1111001101011101", "1111000110100110", "1111101101101110", "1111001110101110", "1110110100010011", "0000010001110110", "1111100111001101", "0001000110000101", "0001001010110001", "1111000010101100", "0001101010100001", "1110001011101110", "0011011000101111", "0000011110000010", "1110101010010110", "1101000010001001", "1110011101100101", "0000110000010010", "0000101111111110", "1111111010101011", "0001110110000100", "1100011000010110", "0000000001010001", "1111111001101001", "0000010000010001", "1101100100001101", "0000001001001110", "0000001100011011", "0010010011000111", "0001010111100011", "1111011001111011", "0000001001000010", "1111001010000100", "1111010110001000", "0000011110101010", "0000000000001111", "1110110001011010", "0000111101110000", "0000110111000111", "0000110000010111", "1111011100010000", "1111110010110111", "0000110111111000", "1111010101011011", "0000101010010001", "1110100110000011", "1110101001111010", "0000110101110101", "1110100110110001", "1111010101111000", "0011101101111100", "0000001111011111", "1110101110011011", "0001100110001011", "1111001100010010", "1100000010110011", "0010101000101111", "0001011010111000", "0011010010101000", "0000111111000111", "1101110010110101", "1100010001010001", "1101000001111011", "1111110101010001", "1110111110011110", "0000011000110111", "0011000011011010", "1110001001001111", "0011010000110101", "0000001011100110", "0000100111110111", "1010101000111000", "1111100000101100", "0000010111111100", "1111101111001001", "0001001000110101", "1110111110001100", "0000001101010011", "1111111011011011", "0001011011110110", "1111101110111000", "1111110010000111", "0001000010101101", "1111101000101110", "0000011011011110", "0000001011001011", "1111111100111101", "1111100110100101", "1110101110101001", "0000110111101110", "1110101000111100", "0010110010111110", "1110100110110001", "0001010100101110", "1110111000001001", "1110100111000100", "1111101101010001", "0000010100100010", "0001100010010010", "0000010101110001", "1110101100001000", "0011100010010000", "0000100111011010", "1100011111111100", "0000011001010101", "1110000111010011", "1111001101101101", "1100110000011010", "1101000001000001", "0001111100110001", "1011110100111101", "0100100010001111", "0100011100010001", "1111001010100011", "0001011100001011", "1111000101110001", "1111101011101101", "1111000110100110", "1111111110110011", "1111111110011001", "1111001011011001", "0000001001101111", "1111011011000101", "1111011111110010", "0000101100011111", "0000011110011110", "0001011100010110", "0000110111001110", "1110011011101001", "0000000100000110", "0000100000011010", "0000000111100101", "1111011011001101", "0000110110101110", "1110000010100011", "0000000111110011", "1101010100011001", "1111101111001110", "1110101110100100", "0100101011001000", "1111011010011000", "0100001000000011", "0001010010100000", "1110011001011001", "0000101100000101", "1101110111011100", "1100001000111101", "0000010100101101", "1111110010110000", "0010011001010110", "1110010000100101", "0000101001100011", "0010001000011110", "1101101011011100", "0010001000011111", "1110011000000011", "1111000000011000", "0000000011000011", "0001110010110111", "0001000101111010", "1111110001101010", "1101110000001011", "0000001011101011", "0000100001010101", "1110110101001111", "0000110100010010", "1110111001101111", "0000011100101110", "1111010110011110", "0000000011101001", "1110010110001100", "0000111001111101", "1110100011110010", "0010111000001110", "1110001010010110", "0000000011111110", "1110010011001000", "1111001011100010", "0000101110101001", "0010001010111011", "1110110101110000", "0000101100101010", "1111011100000100", "0001000101100011", "0000111100001100", "1111111100111001", "1111101100010000", "0000101100000001", "0000011000010001", "1111101101010000", "0000101001110011", "0000101011000111", "0001000100111111", "1111011111101111", "0000000010110101", "0000100111100100", "1111110011101101", "1111011010001100", "0001111100001111", "0001100110100010", "1110111110101110", "1100111111100101", "1101111100010000", "0001010111001010", "1111011010110010", "1111111111110011", "1111101110000100", "0010000001001010", "0010010111101101", "0001011010100101", "1100101111100100", "1110100100001111", "1100000110101111", "0101111110000010", "1111101001110000", "1111101011001010", "0000011100111110", "1101101110111000", "0000100010100101", "1101110011010101", "1101101000110011", "0010100011100011", "1111001100111011", "0010110111110000", "1110111001110100", "1111100000111011", "0000101101101010", "1111000000100101", "1100001001100010", "1111000010000100", "1111011001010111", "0100000011100111", "0001010010110010", "0000010001001000", "1111111001011000", "0000111000010100", "1110100011010000", "1110010100111110", "0001010111011001", "0001101010101110", "0000110101001101", "0001010100011100", "1111100101011010", "0010011000011110", "1111000010101010", "1110100101001111", "1110110111000000", "1111111110100001", "1110101111101010", "1111100000101100", "0001011110000010", "0010001100001001", "1111010001111000", "1111000011011001", "0000001101111101", "0010101011001011", "1110110110001000", "1101101100001000", "1101111101011100", "1111001110001101", "0100100111110100", "1101101010111000", "0001011111000101", "1110001000100111", "0001011101000000", "1111111010101101", "1111101100011110", "1111010010010111", "0101001011000011", "0001010101101101", "0001000000111011", "1111001101111000", "0001101101101001", "0010000111011100", "0000011011100101", "1001111011001001", "1110011000001000", "0010110010010110", "1110111001101000", "0010010010110111", "0001101101111101", "0000110010011100", "1110000100111010", "0001010001101011", "1110001011111010", "0000001000110010", "0000000101110101", "0001011001101100", "0000011001100011", "0000100111101001", "1111101000100100", "0000001100100001", "1111100101101011", "1100000101110001", "1111011110010100", "0000110011100100", "0010001001011001", "1111101011101000", "0000110010001001", "1111101011101111", "1111011001000011", "1111111111111101", "0000010000101111", "1101100000010011", "0000101101100110", "1101101011101011", "1111010111100100", "0001111111001001", "0101001111110110", "1101101011101111", "0010110001010100", "1100100101000101", "1111011111111111", "0000010101001100", "1111001111011101", "1110110110111110", "0000010010101010", "1110111100100011", "0000000101110010", "1111101010100010", "1111110011000010", "1110100101001111", "0000011000111100", "0000000011101001", "1111101110000001", "1111000010001111", "0000010011100111", "1110011011010011", "0001001101111011", "0000100010000100", "0000001101101001", "1110100010101101", "1110011001001111", "0001111110110010", "0001001001000100", "1111111001100011", "0001000000100001", "1111110110101110", "1111111010000101", "0000111010001111", "1101010101010100", "1110111100111001", "1110110101111101", "0001110000000000", "0010010100001011", "0010000000000010", "0001011001000100", "0000110100001101", "1101111100110111", "1111000110101001", "1111100001101111", "0000010010000001", "1111101011000111", "1111010010110000", "1111110111000011", "0000010001111011", "1111001011000011", "0000100011100010", "0010010000011000", "0000100010000100", "1110101010110001", "0000100001111000", "1110101011110001", "0011010001001010", "0000100000000011", "1111011111011100", "1101101110101010", "0001011101110000", "0011111101001010", "0010010111111011", "1101110100111010", "1111111100000110", "1100000001101110", "0010101111101111", "0000110000101011", "1101110010001001", "0001100010110111", "1110000011100010", "0001110010000111", "0001011100011110", "1101010001101101", "0000001100100110", "1111000010100000", "0010101010110001", "1110000110001010", "0000001111101101", "0000001010101011", "1111100010100000", "1111111001101010", "1101111110000110", "1101010011011010", "0011111110101000", "0011001110111100", "0000001011100010", "1110001101011110", "0000000001000001", "1101011100101100", "0000001111010010", "0001011001110010", "0001101101110010", "0010001000110000", "0000111000000100", "1101101111000100", "0010100111110001", "0010001101000100", "1100111110111100", "1010100110110100", "1100100110110011", "1110100110000100", "0001110001101101", "0100001101001111", "0011111111001111", "1010001000000110", "1111011010111010", "1111101111101111", "0100111010011011", "0010001100111101", "1110100011000011", "0000000101100001", "0010001110010000", "0000011000111010", "0001100010010001", "1110110111001011", "0000110000001101", "1110110111001100", "1111100111100100", "0001000110110000", "0000111010010000", "1111111110111000", "0000000110001101", "1110111110011110", "0001101011111100", "0000110010011110", "1111111100010000", "1111010001001110", "1110100000101111", "0000101111111101", "0001110000100100", "0000000111000011", "0000001001011111", "0000110011010011", "0000011101011100", "0000101100101111", "1101111011010011", "0000011010001100", "0000010000001100", "0000100110101101", "1110010001101010", "1110100001010010", "0010001001110100", "1110001001000101", "0001111010111011", "0001101101011011", "1011101110111111", "1111010111101100", "0001101100011011", "0001010111010100", "0100010010100100", "1110011001110111", "1111111101000111", "1110011100000011", "1111000000100000", "0000100010100110", "1111000001100110", "0000011011111011", "1101100101111000", "1111111111101111", "0001010111110011", "0110001010010111", "1101110101010100", "0000011110001010", "1110110110100010", "1111110011111011", "1111110100100111", "1110001000001011", "1101110010110100", "0000110011100101", "1110111011111011", "1110111010100010", "0001001101000011", "0001000101100101", "1111010101001100", "0001001001011001", "0000110111110011", "1111000111111010", "0000000010010111", "0000101010000011", "1111100010110101", "1111101111010100", "0001010101011111", "1111000100010100", "0001000010101111", "0000111011010110", "0000101011000001", "1110111000011010", "1111111101110010", "1111011001010101", "0000100110100011", "0001001010110110", "1111011010100011", "1110101011100100", "1111100111010110", "0000111010011111", "1110101011001110", "1111001101001010", "1110100111010111", "0000110010001101", "0000011010110011", "0000010010010111", "0000000000001000", "1111000111100000", "0000101000101011", "1111111000101101", "0000010110111010", "1111001110110110", "1111011110101001", "0000001001100011", "0000110110001010", "0000111001011110", "0001011000101100", "1111011110011100", "0000010000011111", "0000100001110111", "1111001011010010", "1111101000101010", "1111010001100010", "0000101011110001", "1111011100110001", "0010101000110101", "1110111001010110", "1111011111110001", "0001011000000100", "1111100010100010", "1110111000101010", "1101110001011110", "1111111110001001", "1110101001101111", "0011001101010000", "0000110101111001", "1111110000101000", "1101011111001110", "1111111100101010", "1111110110010101", "1111110100001100", "1110010101100010", "0000111011100110", "1111101000011110", "0000111110001011", "0000111100011011", "0010110110111001", "1110011111011111", "1110111100000100", "0001101110100110", "1111011011100100", "1111100001001001", "1111111000101100", "0000110010001110", "1111001000101011", "0000001111110110", "1111001110000010", "0000001100110011", "1110000100100111", "0000001110000000", "0000000001000101", "0000111101000100", "0000110001101000", "0010100011010101", "1110101010111010", "0001010011111011", "1110000000100001", "0000010000100101", "0000110000101010", "0000100000100111", "0011001001010100", "1100110011100110", "1110011110111001", "1110000011010110", "0010111110110010", "1101001011000110", "0000000010101110", "1111101001000000", "0000011101111100", "1101111001110001", "1111100001101111", "1101001001101111", "0001101001111101", "0010001010010110", "0001101110010101", "1101001001000000", "1111111011011100", "1100110011101101", "0000000111000001", "0000001101100011", "0001001000110011", "1110011000010100", "0010001110101010", "1111111111110011", "1110011101011101", "0001010001010111", "1111110100001011", "0000001110011010", "0000111011101010", "1111110110110110", "1111100011000101", "1111010111000010", "1111011010001111", "1111001010111110", "0000010101110110", "0010110000111010", "1101001010000000", "0000100001000011", "1111010000011111", "0000111011100001", "0001101101110010", "0010010011010111", "1101000111101100", "1101011111000110", "0000101101000011", "1100110001010101", "0000011001001110", "0010000101010110", "1111101000101010", "1111010100011100", "0011000101000100", "0010000000111010", "0000001111011001", "1110011101111110", "0000000101010110", "1110101011111010", "0000110011111000", "0000100110000010", "0000100100101001", "1110111011011000", "1110011101110101", "0000000010010110", "0000000110100111", "1111110111100011", "0000000001011001", "1111111011010110", "0000111010111011", "0000100011000100", "1111001011000011", "0000111011011111", "0000000111110001", "0000001110000101", "1111110000111011", "0000101100111101", "0001010111001010", "1111001001011110", "1111000100101000", "1110111001001101", "1111111001100010", "0000110101010110", "1111011011000010", "0000010101110110", "0000101010011011", "0000001000101100", "0010000011111110", "1111000111011101", "1110110110111101", "0000101101001000", "0001110110000000", "1111101011011000", "1111011001100101", "1101011110010101", "1111110100100101", "1110110110000111", "1111011010111000", "1110101110111011", "1110101111010101", "1111011110000010", "0010110101010011", "0000000011100001", "0000010011010110", "1101110000011111", "0000001001100100", "0000001010100101", "0000100011001100", "0001100111010000", "0000110001010010", "1111000011100110", "0000111101100111", "1111110111001011", "0000011001111100", "0000110111111010", "1111101010001110", "1111110001100101", "0001110001101100", "0001000010101010", "1111100101000000", "0000111111110100", "0000101100001100", "0000011001010111", "0001100011010111", "1101011000100100", "1110010110111001", "1110000110000001", "1101110010001111", "0000011111001101", "0001100011111000", "0000101000110010", "1110110100010011", "1110011000101101", "1111010111110001", "1111110101001100", "0100111110101001", "1110111110011111", "1111010001011100", "1111001001111111", "0010010100110011", "1111100011010001", "0000011101101001", "1111010101100101", "0000001001111011", "0010101101111001", "1111101010110000", "1110100110011101", "0001000011100111", "1111111000100011", "1111000011101110", "0000100011000111", "1111101010001010", "0001001000100101", "0000100000100110", "1110011101011101", "1111000101111100", "1111111001110100", "0000110110111000", "0010011010100011", "1111000000000110", "1111101101001011", "0010010110000010", "1101111001101110", "1111100100100011", "1111010100100000", "0000111110001101", "1111111011111111", "1101101000011110", "0000101001110010", "0011000100110001", "0000101100111100", "0000100001100101", "0001001011011010", "0001000000001011", "1111100011100010", "0010000000110101", "1111111111001110", "1110100011101101", "1110101011101101", "1111000011110100", "1111000100101101", "1111001001001011", "0001010101000101", "0000101101011101", "0000111010101011", "1110011100111001", "1110110010011111", "0000011100101010", "0001000101100110", "1111110000001011", "1111111001101011", "0000101010001011", "0000100001010111", "1111100001011100", "1110110011101010", "0001000010000000", "0001111101000001", "1110101010001101", "0000101101101101", "0000010010010011", "1111010010010010", "1111111110100010", "1110111011010111", "1110001001110001", "0000010011111111", "1110101010011000", "0001011011011101", "1111001111101101", "1111110110011001", "0001000110001010", "1101011011000001", "0001101111011010", "0010101001111110", "1100001100011111", "0011100101001001", "1101100010011000", "1110110001110101", "0001011101010001", "1111010010100001", "0001010100100000", "0000010101010001", "0001011101100000", "0000000001011101", "1101100100000001", "0001001101010001", "1111011101010111", "1110101010101000", "1110111001100001", "0000101100100011", "1111101011010011", "1111101101000101", "1110100011011000", "0000010101000001", "0000111111101001", "1111101010010011", "1111011111011001", "1110111010100100", "0000101110000111", "0001001001101101", "0001100100110100", "1111110000011110", "0000010111011000", "0000100001101011", "1111100111110101", "0000101101101000", "0000010100101010", "1111100101010000", "1110110000010000", "0001100010011100", "0001000101010101", "1111111001111111", "0000100000010100", "1111110001111011", "0000001010000101", "1111011000111100", "0000010100111010", "1111101110110010", "1111011100001001", "1111100110011110", "1110110100100010", "0000011001110110", "1111111000010001", "0000110111011000", "0000110010110010", "1110111010000101", "1111101011010001", "1111010001011101", "0001111000101011", "1101111011000011", "1111101001010010", "0000001110110000", "0000011010100000", "0000000001111111", "0001010000010101", "0000110011110111", "1110010101110100", "1111001111110111", "0010000010100001", "1110110010011001", "1100111110011011", "0001001100100100", "0000110100101010", "1110010000010101", "1111111111100100", "1111000100100000", "0000101110100001", "0100010000010011", "0001011110101000", "0001001111001011", "1111011000100101", "0000100110110000", "0001111010110110", "1100011000110001", "0000000001000011", "1100110100001011", "1110111101000111", "1111110011001110", "0000100011010100", "1111101010101110", "0000100001100111", "1111011111100001", "0000010111111101", "1111111001100101", "1111000100101111", "1110001000100111", "1101110010010010", "1111111001000010", "1101101010010011", "1100110010001001", "1101000100001001", "0010101100010000", "1111100110001110", "1111101010100111", "1101111010111010", "0010011001011111", "0011100000010000", "0000011110100011", "1111111011111101", "1100111100101100", "1110001111110110", "0010000000111001", "0001011000111011", "1110100110101011", "1110110000110100", "0001011100100101", "0010110111001010", "1111101001100101", "0010111110001011", "1100011000010100", "0001011111111000", "1111111001010010", "1110110110110011", "1011011001011000", "1110111101110110", "0001011000101110", "0011000011111011", "0001001110100000", "1110101110010111", "0000010010111111", "1111110111001000", "1111101110010101", "1110100110100000", "0000110111110011", "0000100110011001", "0001001101111011", "1111101010111000", "0000100010101100", "1110110000101001", "0001010011101111", "0001110100101010", "0000010111111111", "1111110000101111", "0000110101001111", "1110011110111001", "0001000101011110", "1111010001110100", "0010000110110011", "1101101110010001", "0101001011110100", "1110111010010011", "0000100001000100", "0000001111011010", "0010001101110110", "1110001110010110", "0001010010011101", "1110000101001110", "1110001101000111", "1111111000101101", "0011101001000100", "1111111000101100", "1110011011001000", "1101110011110000", "0001011010101111", "0000100100111110", "1111000010110110", "1111011011001100", "0000110111110101", "1110100110010100", "1111010010011011", "0001010111111010", "1111100001100001", "0000111010011000", "0001010100100101", "1101001011111111", "1111101110010111", "1111000011111001", "1110111011010101", "1110101110000010", "0010000111001110", "0000110111110011", "1111010010001110", "1110100111010011", "1111100100001100", "0000010111011100", "0000101001110100", "0000101011100100", "0000101001000100", "1110000100001111", "0010111110100110", "1111001100010101", "1110101111110010", "0000011010000100", "0001100110010010", "1110000010101000", "0001000101000001", "0000000001000111", "1111110000000011", "0000111110001000", "1110111111000011", "1110011110111100", "0001010101010101", "0000001111100110", "0001001111011000", "1111100101000000", "0000001101011100", "1110001011100011", "1110111011001101", "0010011100100001", "1111010000011010", "1110100001011010", "0011001100100100", "1110001110110000", "0001011000001001", "1111110000110101", "0000111000010011", "1111010001110001", "1111111110010000", "0001001100000000", "0000011010011010", "0001010111100011", "0000001010011100", "1101110011110111", "1110001100011001", "1110110101110001", "1111100110010010", "0010000011110000", "0001011011100110", "1100101010110100", "0000001100001001", "1110100111101000", "1011111010110001", "0000111111001100", "1101100011011000", "0000010011000111", "0001100010101000", "0011110010000000", "1111001000010101", "0000000011000111", "1111101000001110", "1100000110101001", "0000010100101001", "0000101011010110", "0100000111000010", "1111011110011100", "0001001100111101", "1111101011011100", "1110010001011010", "0001111101011000", "1110111010111000", "0000110101100101", "0101110000010000", "1110111110111010", "1101111000110110", "0000111110110101", "0000000001110011", "1011000001011110", "0000100000101100", "0000001111000011", "0010101100000011", "1111110000111010", "0000110111110100", "0000111001111100", "1110011000011010", "0001111100011010", "0000110111110110", "1101011010100010", "1110110111010110", "1111011111000001", "0001100110010111", "0000010001000111", "1111111001111101", "0000001011110111", "0000010000101000", "0000110010110001", "0000000100011111", "1100100110100110", "0001000001100000", "0010110001010101", "1101101101011101", "0010001001011101", "0001101011010101", "1110011110000011", "0010101001001111", "1101100100100111", "1111111110101100", "1110111111111100", "0001111001101010", "0001111101110110", "0001100110100011", "1111000110011111", "1101111110101111", "1111000101111101", "1101010111110000", "1110010010111000", "1111011001011101", "0011000101010100", "1110000110110011", "0011010011111010", "1111000011010101", "0000010100101111", "0000011110000010", "0011011011010101", "1101010101110001", "1111110110011110", "1101100110100110", "1111010001111110", "1111001010110100", "0000000001101000", "1110111111101001", "1111101100011001", "1100101110100010", "0000001011111001", "1110100100011010", "0010100100100110", "1101111101010100", "0000111000110100", "0000110011010100", "0001000001101111", "0000000001100101", "0001000001101110", "1111001011010000", "0001110101101000", "1101100000000101", "0001001010111101", "0000011010100001", "0001011100101101", "1111011000111110", "0000001000001100", "1110000011011011", "0010011011011111", "1100100101110101", "0010001011100001", "0000010011100001", "0000001000000101", "0010100001011010", "1111110101000110", "0000011001000110", "1111111001010011", "0000100011010101", "0000000011000100", "1110100010100011", "0000101101111100", "0000001110110010", "1111101100111000", "0000111110110101", "0000011111110110", "0000110111111110", "1111010001011010", "0001010110110111", "1101011010101000", "1110110111100101", "0010000011110100", "0000111111111010", "1111100100100001", "0000000011011110", "0000001110111000", "1111111011110000", "0001011101111001", "0000000110011110", "1111100001100001", "0000000011100111", "0001010010101000", "0000011010011101", "1111101111000011", "1110110100110111", "1111101010100111", "0000001100011101", "1111101011010111", "1111011011001010", "1111100000001101", "1111001101010010", "1111011000010001", "0000111111111111", "0000011101001010", "0000101100111010", "0001000010001101", "1111111110011110", "1111001011110100", "0000000001010111", "1111011100000110", "0000110000111011", "0001010000001110", "0000110101001110", "0001001001100101", "1110011010010110", "0001100110101110", "1110000000101100", "0000001001000110", "0000110110110110", "0011111100011000", "1101110110100000", "1111000001111100", "1110111110111111", "0000011010111010", "1101110110000101", "1111001000111100", "0001100101001011", "0001101010101111", "0001100000011110", "1111000101000111", "1101100011101101", "1111000100001100", "1101001101111011", "0100001010100111", "1100001110101110", "1110001000110010", "0001001111001010", "0010000011000101", "0001011100100111", "1101001101001111", "1111010101011000", "1111010101111111", "0001100111101110", "0001010111100111", "1110100101101011", "1110100111000011", "0010001010011010", "1111010110100011", "0000100100011111", "1100011001000101", "0000100010111111", "1111100000010001", "0010001001000010", "1111101110001110", "0000010111000110", "0000001110100000", "1111100100011010", "0010001011010110", "0000111101100001", "1111100101001101", "0000011100100101", "0000000000100100", "1111001101111001", "0000101101110010", "0001111011000110", "1110101010101100", "1110101100010011", "0001011100001000", "1111111011011101", "1111110001100001", "1110111110001001", "0000010011100110", "1111111011111010", "0011010101000001", "1110010110010101", "1110111110001010", "0001000100110011", "1111111110111101", "1101110001010010", "1101101011110000", "1111000001001101", "1110110110101001", "0000111101100100", "1111110101101110", "0000001111001100", "1111101111010000", "0000101011101101", "1111111101000010", "0010001101110100", "1111010000011100", "0000010100110110", "1111011110110011", "0000100010011111", "1100101111011101", "0001011010100000", "1111100110010110", "1100011100111011", "0001000100000110", "1111111110011010", "1011011100101011", "0010110100110110", "1110110001100100", "0000100100111001", "0010101110101000", "1111110111111111", "0000001001101111", "1111000111101010", "1110111000001000", "0000101010000100", "0010100001011101", "0010100010111011", "1111111110110110", "0000010000111000", "1111011010010100", "1110001001010001", "0000101010011011", "0010101001001101", "1111000100000101", "1110111001000001", "0000111100000111", "1111000011010010", "0001111100111011", "0000000101010110", "1110101100100010", "1111001101001000", "1111001011110000", "1111101101110011", "1110011010000110", "0001011110101011", "0000000000010101", "1111111010010111", "1111101000001110", "0001011100100010", "1110010101011101", "1111111010100010", "0000111000010111", "1101011011001000", "1111100011110100", "0010010100111100", "0001100110101001", "1101101000010001", "1111011011000001", "0001100010001100", "1100001000010001", "0010010011010001", "0001000111111101", "0010001111001001", "1111101101010011", "0000101001011000", "1110101000011111", "1111000000010100", "1101110101100101", "0011000111001000", "1101001100101000", "1111001101001010", "0011010001001011", "0001010011111100", "0001111000010000", "1111010101110111", "1110001000011110", "0001111011010011", "0000011010100000", "0010001000110111", "1111001101000001", "1110110100001011", "1110101110100011", "0000010111100001", "0000111100110001", "1110000011011101", "1110111000001001", "0001101010010100", "1110100001100001", "0001010001001100", "0000111111110010", "1111110010011001", "0000011001101010", "0000001010100010", "0000011101101001", "1111011111000011", "1111111000000010", "0001001100000101", "1111001010011010", "1110111111010010", "1110101101011101", "0000001110010110", "1110101000111011", "0001010000110011", "0000111101101010", "1110101011100100", "0010111001101111", "1101110111100000", "1110110111011110", "0000110000110100", "0000100000011010", "1100100110000101", "1111010000010010", "0000100010101011", "0000110101001010", "0010110101010111", "0000000101010010", "1111010110100110", "1111100110000110", "1110011001000011", "0000001010111010", "0001011110001101", "1110101001010100", "0000001011011001", "1111000111110011", "1111011001111010", "1011011001100101", "0010110101001000", "0000111101110001", "0001101001001101", "1111101111100011", "0001000011110011", "1110000110111011", "1111010000011111", "1110111101101110", "0000110111100001", "1100001101100000", "1111100111111100", "1110000010011010", "1111000100110001", "1110100010000010", "0111111111111111", "1110010100010110", "1110111001110001", "1111010100101111", "0011010000001011", "0001010110011000", "0000111010010111", "0000111111001110", "1101001010000110", "0001100010001100", "1110100001010010", "0000100001100100", "0001100110100010", "1111010110001000", "1110011101110110", "1111010100110000", "1111010100010101", "1111111101001010", "1110010100111010", "0000101011110100", "0000000001101001", "0000010010110111", "0000010011010110", "1111000001110001", "0000110101011111", "0000001100000000", "1111000111101011", "0000011110000011", "1111100011100110", "1111111110011001", "1111001101110000", "0000011100111001", "1111010101011011", "1111011011100001", "1101010110111111", "0001101100011111", "1111101110010001", "0001100001111111", "0001000010100001", "0000110110011001", "1110000110110000", "0000110111100010", "1101100000100110", "0001010110111000", "1111011000010100", "0100000101011000", "0000111100010010", "0001011101101110", "1110101000001100", "0001101011101001", "1101100111000110", "0011000010100111", "1111111001011000", "0000100101000110", "1101110110110101", "0001100111010110", "1111100111110110", "0000111111100010", "1111011110000001", "0000100010101011", "1111011110011011", "0000011100101111", "1111101110111011", "1111101000010111", "1111000110110011", "1111111101000001", "0000000110000101", "1111110101010001", "0010000000010000", "1111000111111000", "1111111011111001", "1110000110100101", "1111111101111000", "0001101011110111", "1111001011010001", "1111010100011010", "1111100100000111", "0001011001001101", "0010000110111001", "1110101111100110", "1111111001001001", "1110111011010010", "0000001000110011", "0000111000010001", "0000111110011001", "1110110001001100", "0000111101000001", "0000010100100000", "0001101101011111", "1110100100101100", "0000101100100010", "1110000000000010", "1111100010100110", "0000011000101000", "1111110001100000", "0000010010011010", "1111100100010110", "0000010100011010", "0001100011001010", "1111010011110100", "0000110000110100", "1111010110101010", "0001000000101011", "1111001000001010", "1101101001101111", "1111011011110101", "1111000111100001", "0010100110011010", "0000111000000011", "1111101010011111", "0001011110100010", "1111010011000001", "1111100101110001", "0000101110111010", "1111011010100100", "1111001000111010", "0001101100111010", "0001101111010010", "0000101011101101", "1110000100010010", "0000000111111101", "0001001010101110", "0010000001011100", "1111010001011101", "0001001101010100", "1111101001001110", "0001000100110101", "1110111110100111", "1110011011101011", "0010100111100000", "1101000010000100", "1101000111010110", "0001010011111010", "1110011010101001", "1110010010000010", "0001101001101011", "1110111101110010", "1111100111011000", "0000111100110010", "1111111011011100", "0000100010011100", "1110001000001100", "0000000010000110", "1101001101100100", "1101100010011111", "1110111111010001", "1111110111000110", "1111101010100101", "0011001110001010", "1110100101010110", "0010000111011101", "0001011010111001", "0000010011010101", "1111101010000101", "1110001001010110", "0000011110010011", "1110110000000111", "0000000110010000", "0000101101110111", "1110100101100111", "0000011100001110", "1110101100101011", "0000101100010111", "0011010000100010", "1101101000010100", "1110000000000111", "0001001010100011", "0001000010001101", "1100101001000111", "0000011011111100", "1110110001010011", "0001110011010000", "0000101010100101", "1110101100110111", "1111010001101101", "0000011000010000", "0000111111101110", "1111110100110011", "1111010001100011", "1110110100110111", "1111001101010100", "0001011110000010", "0000100110011001", "1110000000101111", "0010001010110000", "1111101111100001", "0001000100001110", "1111100001000011", "0000100110111011", "1110100111000111", "0001011100100010", "1101100011101110", "0000110111001100", "0000000011111111", "0000101100100100", "1101110000011111", "1110110110110110", "1011111001011011", "0001110011011011", "0001000000101010", "0010001011000110", "1111101010000111", "1010000001010001", "0000011000110010", "0001010111101110", "1101111011100111", "0110001011100111", "1100110011110111", "1100111100010000", "0100101000110010", "1101111101001111", "0101101011111001", "1101111111010111", "1111010110010111", "0001000001000101", "1111100000110100", "0001110111011100", "0000001110101000", "1111001111101100", "1111000101001011", "0000010001001101", "0001100001110110", "1111011100100010", "1111100110110101", "1111011100111100", "1111100101011110", "1110100101110000", "1110100000111101", "1111010010101111", "0001010001011100", "0000010010111011", "0000101010010000", "0000010110110100", "1111110010100011", "1111011011110101", "0000110111011000", "0000000100001100", "1110100111111110", "0001010010010101", "1111010111010100", "0000011010110001", "0001110100110101", "1101100011100101", "0000110111001100", "0000011100000111", "0011010010001110", "0000000110100011", "1110100001010100", "0000110011101000", "0000001111001111", "1110001101110010", "1111001001010111", "1101101101010101", "0000000001011001", "1111110110011010", "0000001110010001", "1111110001100100", "0001011010101000", "1111111111011011", "1110101001010100", "0000010111010111", "1110111111011000", "1111001110010100", "1111001001010010", "0000100000100111", "1111100110110100", "1110111011101001", "1110111110101100", "0000001100010001", "0000001011001001", "0000100111111000", "1110101010110101", "0001110010101010", "0001100000001011", "1111000001111100", "0000011110101000", "1110111111100000", "1110001000100001", "1111011010100001", "0000000000100000", "1111111000001110", "1110011010011000", "1110011111001001", "0001000101101110", "0001101100010100", "1111110100101110", "1111110111011010", "0001000101011110", "0000110011011000", "0011101000110100", "1110101100001100", "1110001010110101", "0000001000111101", "1110010010110000", "1111001110000101", "0001100111011010", "0010000101101000", "0001101110001110", "0001001001111110", "0000000010101111", "0000111110100110", "1111000000011000", "0000001000001011", "1110111110100110", "0000101011100011", "1110001101010111", "0000101011100100", "1111101001000101", "1111101010111010", "1111111011101000", "1111001000110111", "1111000101100010", "1110101110100111", "0001110010000110", "1111000100110110", "1110100111100010", "1111110110011011", "1111110111110110", "0000000110011100", "0000001100100000", "0001001011111111", "0001010101010111", "1110010011110001", "0000000111100001", "1110011100110010", "1110110001110101", "0001010111010111", "0000100110010000", "1111000011000101", "1111001101001101", "0000010010101100", "0010011111010000", "1111001110111001", "1111001011110000", "0011100110000100", "1110011100110101", "0001111010010000", "1110111101111011", "0000001101110000", "0010000011011000", "1110011010010000", "1110111110001011", "1111101111111000", "1111001001100110", "1111101100100000", "0000010000011010", "1111100000000101", "1111010110101111", "0001000100001100", "0000101010010111", "0000101010000101", "0000001111111011", "0000000101011110", "0000001111011101", "1100010011100001", "0001011110000010", "0000001011000101", "1111010111000001", "0000001000101100", "1111101001010110", "0000100110110100", "0001000110110111", "0001110111110111", "1111110101110011", "0000100010011110", "1111011100010011", "0000011001110011", "0000010011011110", "1111000001011101", "1111010011011000", "1111011111011000", "0001010110111010", "1111000111011110", "0000011110001110", "0011101011000000", "1110110110010011", "0001001101111000", "0001001010000101", "1111011000111011", "1101100101110111", "1111100100111101", "0001110110000010", "1110001101001110", "1111001000011100", "1111100111110011", "0001000110101001", "1101111110110100", "0001001110110010", "1111010110001111", "0001011011011001", "0001111000110011", "1110100011110000", "0000011100110110", "0001011101010011", "1111100000111011", "0000010010000110", "1111010101000101", "1111111011000000", "1111001001110101", "1111001100011110", "0000100101110011", "0001010011001100", "0001010011001110", "0000100101001100", "1101110111000100", "0000100010010011", "0001100100001010", "0001011001000100", "1101010101111111", "1110010011010001", "0000001011000000", "1111101011010011", "0000101010011010", "1111100110100101", "1111101010010111", "1111100100100100", "0001111000001001", "0010001101000000", "0000010011001010", "0001111001110100", "0000000111100001", "1111001011110111", "0000101011011000", "1111100101110100", "0000001101000011", "1100110011001111", "0010110000000101", "1111011001111110", "0000110010010011", "0001001110110101", "1110001010011000", "0001011110111001", "0000011100010100", "1111110001111000", "1111001111110110", "1111000111011011", "1111010101011000", "0001010100110010", "0001100010101110", "1110101101000010", "1101101110010010", "1111111110001111", "1111001000000001", "0010000111111010", "1111101111000010", "1111010000001111", "1110111000111011", "0000100100010010", "0010000101000011", "0001011000001110", "1101111101011100", "1111100010111111", "0000100101011100", "1111100001010110", "1111010000111000", "1110001100100110", "1110110000111011", "1111111111011010", "0010001000101010", "0001000000100010", "0010100100111111", "1110111101110001", "0000010101000001", "1110110001101111", "0011101111011001", "1101111111101110", "1111010110101010", "1110110011111111", "0000100101110100", "1101011001001111", "1111011101011011", "0000000011111100", "1111110111111101", "0001111001000011", "0011101101000110", "1101110001001111", "1110110011100101", "1111011000101101", "0001111000101010", "1111100101100111", "0100000001001001", "1011110101011011", "0000000100110000", "1111111010011111", "0011000100100101", "1110101111001011", "0000001101101101", "1101111111100110", "0001000100011101", "0000000111001110", "1110001011001110", "0011000010111111", "0000101010001011", "1111100110001111", "1101110000110111", "0001001100110010", "1110111101111101", "0000110100001100", "1111010010010101", "1111010111000010", "0000000011100001", "1110110101110101", "1111000011011101", "0000101100010000", "1111000000110110", "0011000111111010", "0000000001100100", "1111100110100011", "1110001111111111", "0001001110011001", "0001000100100011", "0000111011000111", "1111101111100100", "1111001010001111", "0001101011010110", "1111110001010000", "1110001100001100", "0000110001100011", "1110001111001000", "0000111110111101", "1110111000110010", "0000010110000000", "1111001101010110", "0000100001011011", "0000001111000000", "0000101011111101", "1110011010111111", "0000110010001000", "1111110010001001", "1110110011110010", "1111110011000010", "0001111010011011", "1111111001000110", "1111001100111110", "1111010001010101", "0000001000001110", "0010001101111100", "1111001010001100", "1111001110111010", "0000010101101100", "1111100110000111", "1110010011001000", "0000111100010001", "0000011011001010", "1110110100010001", "1111110010010011", "0000101111110011", "1111001100000011", "1111110011100110", "0000011001101110", "1111111011000100", "0000110110010000", "0000101001001010", "1110110011011100", "0000100100111010", "0000101010000110", "1111010000010111", "0000101111101111", "1101110000111110", "1111111011000000", "0001010011001111", "0000010111010000", "1111111110111111", "1111011100101111", "1110100000110010", "0000000010010110", "1110010110000001", "0000011101000101", "0001010011011100", "1110101111010011", "1111001100110000", "0000100011000000", "1111010101000110", "0000011111110000", "1101111010011110", "1110100010011010", "1110110000110101", "0001110001010111", "0010011000011010", "0001001000101110", "0000001101110100", "1110011111011111", "1111001010101011", "0000111001010010", "0001100010100110", "0000111101111101", "0000000001111111", "1111101010100111", "1110111110011010", "0000000011001111", "1111000000011000", "1111100100011111", "1111100001100011", "0000010001010101", "0010001100001000", "1111111100100011", "1111001101110000", "1111110000010100", "0000110011110111", "0000100011010111", "1111110101000111", "1110010110000111", "0001010010000101", "0100000010011111", "0000111111111100", "1111000101000001", "1110001100100010", "1111111000101001", "0000101110101010", "1110110000100001", "1110010100111010", "1111001111001100", "1101011110010110", "0001010000110011", "1110111001100100", "0000111000100000", "0000000000011001", "0001011001101110", "0010010011001010", "0001010010100111", "1110100000010000", "1111010100011100", "1101111101011100", "0000110011011100", "1111010010100011", "0000001000011110", "1111011110101011", "0001000110001110", "1101111110110010", "0001111011111010", "0001101010010000", "1111101001101000", "0010000100011000", "0001011010110101", "0001000100111100", "1101011100011110", "1111110011001111", "1110000001010111", "1110001011000011", "0010010110010011", "1110101110111011", "1111111101101100", "0000100100111000", "0010100100101100", "0000100100100000", "1111111110110101", "1111001001001110", "0001010110011000", "1111111111100010", "0010001010011110", "1111001001010000", "1101110110000010", "1111010000001100", "1101001010110100", "1101100101111011", "0010110100010101", "1111011110000011", "1101011101011011", "1110001011011010", "1111100011101111", "0011110011111000", "0010100001010010", "0000000011101111", "1100111010011100", "1111001100011101", "0001001100100001", "0000001111111011", "0000101011101110", "0000101101111111", "1111110011000011", "1111001101110110", "0010000101101010", "0001100100111010", "1111111100000101", "0011111100111110", "1110100010010000", "0000111000111111", "1111010001110010", "0001010101110101", "1110001000100101", "1110010000000000", "1110011010101011", "0000111110010010", "0000100010110000", "0001001010000100", "1110001111010101", "1111101000001101", "1111110101011010", "0000000000101001", "0001001000110001", "1101111111100011", "0000000111111010", "0010110000101111", "1101001110101011", "0000001010101100", "0010011101111100", "0000011110000001", "0000010111110110", "0001110001010110", "1111000000011111", "1111011000001110", "1111011001101110", "1111001001000010", "1111011001111000", "1111101100101011", "0000100000110000", "0000111010000011", "1110111001100110", "0001010101001110", "0000010000101010", "0000110111000110", "1111101011000110", "1111111110101111", "0010011101000110", "1110101001110100", "1101101110100101", "0010110110111101", "0001001111100101", "0001011101011111", "0001001010110110", "1110100011101100", "1110000011000100", "1111011101100001", "0001001010111101", "1111110000000000", "1100111110000001", "0010111010101111", "0000101101001010", "1111011010110111", "1111011100000100", "0000000011111110", "1100100100011011", "1111010000111001", "0011001000100011", "1101100000011111", "1111000101001001", "0001111010100011", "0000101001110001", "0000101111001110", "1111010110111011", "1111011101010001", "1101011011011010", "0001101100010001", "1110111011101101", "1110000111101010", "1110100100010000", "0000011111001010", "1111101010000011", "0001101111001011", "1110010110011010", "0001100110111100", "0000101001010110", "0001110010101111", "1011010111101111", "1111100111011000", "1110000110110100", "0010101100101010", "0001001001000010", "0010011000000010", "1101110110000001", "0000011001111111", "1111111000010110", "1110111010100100", "0000001000000001", "0000000111001100", "0100010100100111", "1100100110001111", "1101111011010001", "0000011101101010", "0010000110111111", "0000101001001001", "1110000011101100", "0000111101110000", "0000101110000001", "0011111010100001", "0001011011101110", "1111100001000011", "1010100010100111", "1101111001001110", "1110111001010000", "0010001111011010", "0001000101101001", "0010001110101001", "1110110110111011", "1101000101011001", "0000000101011101", "1111101000001111", "1111000110100101", "0001110110000100", "1111011100000011", "0010000000101000", "0000111100110000", "0010010100001101", "1101011111010110", "0000111001100101", "1011110111100110", "0010110111000001", "1110011101000110", "1110100101100110", "1111100111011111", "0001001111011111", "0010111011101110", "1111001101100110", "1111101000000100", "0001100100010101", "1110111011101010", "1111100100000110", "1111111011101000", "1110010111001011", "1110010111000100", "1110100111010001", "0000010001000011", "1111100001111011", "1111111101100001", "1110011110110111", "0000111100110011", "1111010001011111", "0000110000010000", "0001001000011011", "0001110001000100", "0000001110001001", "1111100011001111", "0001010001001101", "1110110110000101", "0001010100001100", "1110110001101100", "1110101010011110", "0000010101011101", "1111010000111010", "0000110000111111", "1111110010100001", "1111101001011001", "1110100110101111", "0010010001100000", "1100000111100000", "1101101001011001", "0010000110011010", "1111010010111000", "1110010010110010", "0011100010110001", "1111001100100000", "0011001001111011", "1011100101110101", "0000011110100000", "1110110001100001", "0001000100010100", "0011110010001011", "0000010111011000", "1110011110111010", "0100010111110001", "1101001101001101", "0100000001011111", "1101110111111001", "1111010111011001", "1100111010110110", "0010011100110101", "0001010101011101", "0000110010100111", "1111111011010011", "0000011100100110", "0001110011011011", "0000010010000011", "1111100100000100", "1111111101011110", "1110111100001111", "1111001011110010", "0000001111111011", "1111110000100000", "1111010100101111", "1111101100100101", "1111001010110011", "1111001110011100", "1111001100000111", "0010100101101111", "1101110110011110", "0000011001011110", "0000110110011001", "0000000010101010", "1110101101000101", "0000110011100011", "1111100100010101", "1110010100010100", "0000111101001100", "0010000110000001", "1110111010011111", "0000000100000101", "0010111010101000", "1101101011010000", "0001001101011011", "0000001111110100", "0000101110100100", "1100010011000010", "1110010000100010", "1111111101011001", "0001001010100011", "0001101101110010", "0001101001011111", "1110110111101101", "0001010000111110", "1111111011100011", "1111001101110010", "0000101000101100", "1110111000100000", "0000011111100110", "0000100010010110", "1111110111010111", "0000110010100110", "1111100011011001", "0000000111110111", "0001000101011100", "1110111111111101", "1111101111011010", "0000100010111000", "0000011010011000", "1111010010001001", "1110011100111110", "0000010100100011", "0001000000100100", "1111110101010011", "0000010011100111", "1101110110100110", "1110101010001001", "0001000100001100", "0001100011111110", "1111110010001001", "1111111001000000", "0001001100010101", "1111000111100100", "1101110111000000", "0001010111010100", "1101100001000111", "1110111101010010", "0000011001001111", "1110101110100011", "1111111000000001", "0000011010001110", "0001000111100100", "1111001010000100", "1110110100010101", "1110101001100111", "1111011000101111", "0010000000010000", "1111111110011110", "1110100100111000", "0000000110010000", "1111100010100100", "1111000111011111", "1111110010110110", "0000100100111001", "0001000001111101", "1111001000111011", "1111101100101011", "1110110111001110", "1111111000101011", "1111000110100000", "0010111110110000", "1110010101000001", "0001000111010100", "1111001000010010", "0001101001101101", "1110111010001001", "1111110101101110", "0000011011100010", "0000111010110011", "1111100001101000", "1101101101010000", "1110011010111111", "0010000100101110", "1111101000111111", "0001000010000010", "1111101111000110", "0000110101010000", "1111001010010010", "1101000110111101", "1100101111001011", "0100010000110101", "1100011101111001", "0011110010001110", "0001110110010111", "1101010011110010", "0011001111000100", "1110101111000011", "1111001110001110", "1111100011000010", "1111010100110100", "1111011011011011", "0001001111111101", "0001011100111100", "1110101010011011", "1111001111100110", "1111000010001010", "0000001001101001", "0001010011010001", "1111011101010010", "0000011101111111", "1111101001111110", "0001001000111101", "1110101101000000", "1110100000111101", "0000011110100101", "0010001001001000", "1111110001110010", "1110111100101010", "0001011001101010", "1110110010110110", "0001000010110101", "1110101000101011", "0000100111111001", "1101101101111110", "0000111110100100", "1111010000100101", "0001000110010000", "1110011000000101", "0000000001110011", "0001100000010001", "0000001110100101", "1111111011001100", "0000001011100111", "1111001101101100", "1110100011100100", "0011101111011110", "1110101100110110", "0000110011100011", "1111110110000000", "1111011011101101", "1111101010011100", "0000000011110010", "1111100100111100", "1111000100101101", "1110111111011000", "0000011110101011", "1110110110101011", "1111001010100010", "0000010101001000", "0000111011111110", "1111000010100010", "0001011010001000", "1110100110010000", "0010000011111101", "0001010110000101", "1111110110001100", "1110011101100001", "1110110100010111", "0001001011100001", "1110000110110100", "0000110111011001", "0000011011000010", "1101111110000011", "0011001001110111", "1111111100001101", "1111000010001100", "1110111001000000", "1111001110000001", "0000011000111000", "1110100111110111", "0000011011011110", "0000100010010010", "0000001011010110", "1111111111110111", "1111101111100110", "1111100001100000", "0000100010001000", "0000010011011001", "1111011011001000", "1111111000100101", "1111001101010101", "1111100010001101", "1111011100011001", "1111100000000001", "1111000111111100", "0001000101111001", "0000110110011110", "1110101000111111", "1110011101100111", "1101100000101110", "1111011101110111", "0010001001010010", "1110100000101110", "0011001011100110", "0000001011111100", "0000011101100001", "0001101111001111", "0010000101100101", "0000100010000110", "0000000010100110", "1011111010000011", "1111101101011101", "0001000010101001", "0010001110010111", "0000010000100001", "1101000000111101", "0000000110011100", "1101101011110110", "0010000111010101", "1110011110000010", "0000100000110011", "0011011111110101", "1100111111011111", "1111000011101000", "0010001010111101", "0000101000001000", "1111001001101001", "0000011101010100", "1111110011001010", "1111101111010110", "1111001101100110", "1111101010000011", "0000100010010001", "0000001001110111", "0001000010010010", "1110111100101101", "0000110100000000", "0011001010001001", "1110001111011110", "1101010110110000", "1101111011001010", "1111110010110101", "1110011111111011", "0000010100100100", "0100001001000010", "1111101111011110", "0000010000111100", "1111011110000100", "0010111101001101", "0000101100001110", "1110010000101101", "1101011000010011", "0001101000001000", "0000010101010100", "1111101100111010", "0010000011010001", "1101111010010110", "0010011000010101", "1110111100001001", "0010110010100010", "1100110011001011", "1111110011110011", "0001001110010001", "1101001100100000", "0011001101100100", "1111111101000111", "1101111101000010", "1111110000010001", "1111000001111000", "1110110111100110", "0000011110010000", "1111010011010111", "0000101110011000", "0000000100101001", "0000000011010101", "0000000011000010", "1111111011101111", "1110100100111100", "0011100110011001", "1110110000100001", "1110010100000111", "0000100010000110", "0001010011000111", "1111011110101100", "0000000000101101", "1110100001011000", "1111000110010001", "1111001100100001", "0000110010010000", "1110011001011100", "0000000010110110", "0010111010010011", "0000111001100110", "1100010010101001", "0000011111011100", "1101000000101011", "0100001001101001", "0001000001111100", "1111000011011111", "1110111000110101", "0001101010011001", "1101110100101101", "0010001010001011", "1110001110011011", "0001111000010111", "1111101101010010", "0000111110011110");
    Plus214_i_1 <= ("1111101001000011", "0000000011111111", "0000100010110111", "0000001111010110", "1110111111010010", "0001000111110010", "1111100011101101", "1111100110101110", "0000101011001011", "1111100100000101");
    process(all)
    begin
        next_feedback <= feedback;
        next_state <= state;
		next_was_valid <= was_valid;
        valid_out <= '0';
        output <= (others => (others => '0'));

        case state is
            when 0 =>
                next_state <= 0;
                if valid_in then
                    next_state <= 1;
                end if;
            when 1 =>
                Block386_i_0 <= input(783 downto 0);
                next_feedback(783 downto 0) <= Block386_o;
                next_state <= state + 1;
            when 2 =>
                Convolution28_i_0 <= feedback(783 downto 0);
                next_feedback(6271 downto 0) <= Convolution28_o;
                next_state <= state + 1;
            when 3 =>
                Plus30_i_0 <= feedback(6271 downto 0);
                next_feedback(6271 downto 0) <= Plus30_o;
                next_state <= state + 1;
            when 4 =>
                ReLU32_i_0 <= feedback(6271 downto 0);
                next_feedback(6271 downto 0) <= ReLU32_o;
                next_state <= state + 1;
            when 5 =>
                Pooling66_i_0 <= feedback(6271 downto 0);
                next_feedback(1567 downto 0) <= Pooling66_o;
                next_state <= state + 1;
            when 6 =>
                Convolution110_i_0 <= feedback(1567 downto 0);
                next_feedback(3135 downto 0) <= Convolution110_o;
                next_state <= state + 1;
            when 7 =>
                Plus112_i_0 <= feedback(3135 downto 0);
                next_feedback(3135 downto 0) <= Plus112_o;
                next_state <= state + 1;
            when 8 =>
                ReLU114_i_0 <= feedback(3135 downto 0);
                next_feedback(3135 downto 0) <= ReLU114_o;
                next_state <= state + 1;
            when 9 =>
                Pooling160_i_0 <= feedback(3135 downto 0);
                next_feedback(255 downto 0) <= Pooling160_o;
                next_state <= state + 1;
            when 10 =>
                Times212_i_0 <= feedback(255 downto 0);
                next_feedback(9 downto 0) <= Times212_o;
                next_state <= state + 1;
            when 11 =>
                Plus214_i_0 <= feedback(9 downto 0);
                output(9 downto 0) <= Plus214_o;
                if valid_in then
                    valid_out <= '0';
                    was_valid <= '1';
                elsif was_valid then
                    was_valid <= '0';
                    next_state <= 0;
                end if;
        end case;
    end process;

    process(clk, rst)
    begin
        if rising_edge(clk) then
            if rst = '1' then
                feedback <= (others => (others => '0'));
                state <= 0;
                was_valid <= '0';
            else
                feedback <= next_feedback;
                state <= next_state;
                was_valid <= next_was_valid;
            end if;
        end if;
    end process;
end Behavioral;

